module mult_64x64_lut6_akak(in0, in1, out);

input  [63:0]  in0;
input  [63:0]  in1;
output  [127:0]  out;

wire [5:0]  pp0;
wire [5:0]  pp1;
wire [5:0]  pp2;
wire [5:0]  pp3;
wire [5:0]  pp4;
wire [5:0]  pp5;
wire [5:0]  pp6;
wire [5:0]  pp7;
wire [5:0]  pp8;
wire [5:0]  pp9;
wire [5:0]  pp10;
wire [5:0]  pp11;
wire [5:0]  pp12;
wire [5:0]  pp13;
wire [5:0]  pp14;
wire [5:0]  pp15;
wire [5:0]  pp16;
wire [5:0]  pp17;
wire [5:0]  pp18;
wire [5:0]  pp19;
wire [5:0]  pp20;
wire [5:0]  pp21;
wire [5:0]  pp22;
wire [5:0]  pp23;
wire [5:0]  pp24;
wire [5:0]  pp25;
wire [5:0]  pp26;
wire [5:0]  pp27;
wire [5:0]  pp28;
wire [5:0]  pp29;
wire [5:0]  pp30;
wire [5:0]  pp31;
wire [5:0]  pp32;
wire [5:0]  pp33;
wire [5:0]  pp34;
wire [5:0]  pp35;
wire [5:0]  pp36;
wire [5:0]  pp37;
wire [5:0]  pp38;
wire [5:0]  pp39;
wire [5:0]  pp40;
wire [5:0]  pp41;
wire [5:0]  pp42;
wire [5:0]  pp43;
wire [5:0]  pp44;
wire [5:0]  pp45;
wire [5:0]  pp46;
wire [5:0]  pp47;
wire [5:0]  pp48;
wire [5:0]  pp49;
wire [5:0]  pp50;
wire [5:0]  pp51;
wire [5:0]  pp52;
wire [5:0]  pp53;
wire [5:0]  pp54;
wire [5:0]  pp55;
wire [5:0]  pp56;
wire [5:0]  pp57;
wire [5:0]  pp58;
wire [5:0]  pp59;
wire [5:0]  pp60;
wire [5:0]  pp61;
wire [5:0]  pp62;
wire [5:0]  pp63;
wire [5:0]  pp64;
wire [5:0]  pp65;
wire [5:0]  pp66;
wire [5:0]  pp67;
wire [5:0]  pp68;
wire [5:0]  pp69;
wire [5:0]  pp70;
wire [5:0]  pp71;
wire [5:0]  pp72;
wire [5:0]  pp73;
wire [5:0]  pp74;
wire [5:0]  pp75;
wire [5:0]  pp76;
wire [5:0]  pp77;
wire [5:0]  pp78;
wire [5:0]  pp79;
wire [5:0]  pp80;
wire [5:0]  pp81;
wire [5:0]  pp82;
wire [5:0]  pp83;
wire [5:0]  pp84;
wire [5:0]  pp85;
wire [5:0]  pp86;
wire [5:0]  pp87;
wire [5:0]  pp88;
wire [5:0]  pp89;
wire [5:0]  pp90;
wire [5:0]  pp91;
wire [5:0]  pp92;
wire [5:0]  pp93;
wire [5:0]  pp94;
wire [5:0]  pp95;
wire [5:0]  pp96;
wire [5:0]  pp97;
wire [5:0]  pp98;
wire [5:0]  pp99;
wire [5:0]  pp100;
wire [5:0]  pp101;
wire [5:0]  pp102;
wire [5:0]  pp103;
wire [5:0]  pp104;
wire [5:0]  pp105;
wire [5:0]  pp106;
wire [5:0]  pp107;
wire [5:0]  pp108;
wire [5:0]  pp109;
wire [5:0]  pp110;
wire [5:0]  pp111;
wire [5:0]  pp112;
wire [5:0]  pp113;
wire [5:0]  pp114;
wire [5:0]  pp115;
wire [5:0]  pp116;
wire [5:0]  pp117;
wire [5:0]  pp118;
wire [5:0]  pp119;
wire [5:0]  pp120;
wire [5:0]  pp121;
wire [5:0]  pp122;
wire [5:0]  pp123;
wire [5:0]  pp124;
wire [5:0]  pp125;
wire [5:0]  pp126;
wire [5:0]  pp127;
wire [5:0]  pp128;
wire [5:0]  pp129;
wire [5:0]  pp130;
wire [5:0]  pp131;
wire [5:0]  pp132;
wire [5:0]  pp133;
wire [5:0]  pp134;
wire [5:0]  pp135;
wire [5:0]  pp136;
wire [5:0]  pp137;
wire [5:0]  pp138;
wire [5:0]  pp139;
wire [5:0]  pp140;
wire [5:0]  pp141;
wire [5:0]  pp142;
wire [5:0]  pp143;
wire [5:0]  pp144;
wire [5:0]  pp145;
wire [5:0]  pp146;
wire [5:0]  pp147;
wire [5:0]  pp148;
wire [5:0]  pp149;
wire [5:0]  pp150;
wire [5:0]  pp151;
wire [5:0]  pp152;
wire [5:0]  pp153;
wire [5:0]  pp154;
wire [5:0]  pp155;
wire [5:0]  pp156;
wire [5:0]  pp157;
wire [5:0]  pp158;
wire [5:0]  pp159;
wire [5:0]  pp160;
wire [5:0]  pp161;
wire [5:0]  pp162;
wire [5:0]  pp163;
wire [5:0]  pp164;
wire [5:0]  pp165;
wire [5:0]  pp166;
wire [5:0]  pp167;
wire [5:0]  pp168;
wire [5:0]  pp169;
wire [5:0]  pp170;
wire [5:0]  pp171;
wire [5:0]  pp172;
wire [5:0]  pp173;
wire [5:0]  pp174;
wire [5:0]  pp175;
wire [5:0]  pp176;
wire [5:0]  pp177;
wire [5:0]  pp178;
wire [5:0]  pp179;
wire [5:0]  pp180;
wire [5:0]  pp181;
wire [5:0]  pp182;
wire [5:0]  pp183;
wire [5:0]  pp184;
wire [5:0]  pp185;
wire [5:0]  pp186;
wire [5:0]  pp187;
wire [5:0]  pp188;
wire [5:0]  pp189;
wire [5:0]  pp190;
wire [5:0]  pp191;
wire [5:0]  pp192;
wire [5:0]  pp193;
wire [5:0]  pp194;
wire [5:0]  pp195;
wire [5:0]  pp196;
wire [5:0]  pp197;
wire [5:0]  pp198;
wire [5:0]  pp199;
wire [5:0]  pp200;
wire [5:0]  pp201;
wire [5:0]  pp202;
wire [5:0]  pp203;
wire [5:0]  pp204;
wire [5:0]  pp205;
wire [5:0]  pp206;
wire [5:0]  pp207;
wire [5:0]  pp208;
wire [5:0]  pp209;
wire [5:0]  pp210;
wire [5:0]  pp211;
wire [5:0]  pp212;
wire [5:0]  pp213;
wire [5:0]  pp214;
wire [5:0]  pp215;
wire [5:0]  pp216;
wire [5:0]  pp217;
wire [5:0]  pp218;
wire [5:0]  pp219;
wire [5:0]  pp220;
wire [5:0]  pp221;
wire [5:0]  pp222;
wire [5:0]  pp223;
wire [5:0]  pp224;
wire [5:0]  pp225;
wire [5:0]  pp226;
wire [5:0]  pp227;
wire [5:0]  pp228;
wire [5:0]  pp229;
wire [5:0]  pp230;
wire [5:0]  pp231;
wire [5:0]  pp232;
wire [5:0]  pp233;
wire [5:0]  pp234;
wire [5:0]  pp235;
wire [5:0]  pp236;
wire [5:0]  pp237;
wire [5:0]  pp238;
wire [5:0]  pp239;
wire [5:0]  pp240;
wire [5:0]  pp241;
wire [5:0]  pp242;
wire [5:0]  pp243;
wire [5:0]  pp244;
wire [5:0]  pp245;
wire [5:0]  pp246;
wire [5:0]  pp247;
wire [5:0]  pp248;
wire [5:0]  pp249;
wire [5:0]  pp250;
wire [5:0]  pp251;
wire [5:0]  pp252;
wire [5:0]  pp253;
wire [5:0]  pp254;
wire [5:0]  pp255;
wire [5:0]  pp256;
wire [5:0]  pp257;
wire [5:0]  pp258;
wire [5:0]  pp259;
wire [5:0]  pp260;
wire [5:0]  pp261;
wire [5:0]  pp262;
wire [5:0]  pp263;
wire [5:0]  pp264;
wire [5:0]  pp265;
wire [5:0]  pp266;
wire [5:0]  pp267;
wire [5:0]  pp268;
wire [5:0]  pp269;
wire [5:0]  pp270;
wire [5:0]  pp271;
wire [5:0]  pp272;
wire [5:0]  pp273;
wire [5:0]  pp274;
wire [5:0]  pp275;
wire [5:0]  pp276;
wire [5:0]  pp277;
wire [5:0]  pp278;
wire [5:0]  pp279;
wire [5:0]  pp280;
wire [5:0]  pp281;
wire [5:0]  pp282;
wire [5:0]  pp283;
wire [5:0]  pp284;
wire [5:0]  pp285;
wire [5:0]  pp286;
wire [5:0]  pp287;
wire [5:0]  pp288;
wire [5:0]  pp289;
wire [5:0]  pp290;
wire [5:0]  pp291;
wire [5:0]  pp292;
wire [5:0]  pp293;
wire [5:0]  pp294;
wire [5:0]  pp295;
wire [5:0]  pp296;
wire [5:0]  pp297;
wire [5:0]  pp298;
wire [5:0]  pp299;
wire [5:0]  pp300;
wire [5:0]  pp301;
wire [5:0]  pp302;
wire [5:0]  pp303;
wire [5:0]  pp304;
wire [5:0]  pp305;
wire [5:0]  pp306;
wire [5:0]  pp307;
wire [5:0]  pp308;
wire [5:0]  pp309;
wire [5:0]  pp310;
wire [5:0]  pp311;
wire [5:0]  pp312;
wire [5:0]  pp313;
wire [5:0]  pp314;
wire [5:0]  pp315;
wire [5:0]  pp316;
wire [5:0]  pp317;
wire [5:0]  pp318;
wire [5:0]  pp319;
wire [5:0]  pp320;
wire [5:0]  pp321;
wire [5:0]  pp322;
wire [5:0]  pp323;
wire [5:0]  pp324;
wire [5:0]  pp325;
wire [5:0]  pp326;
wire [5:0]  pp327;
wire [5:0]  pp328;
wire [5:0]  pp329;
wire [5:0]  pp330;
wire [5:0]  pp331;
wire [5:0]  pp332;
wire [5:0]  pp333;
wire [5:0]  pp334;
wire [5:0]  pp335;
wire [5:0]  pp336;
wire [5:0]  pp337;
wire [5:0]  pp338;
wire [5:0]  pp339;
wire [5:0]  pp340;
wire [5:0]  pp341;
wire [5:0]  pp342;
wire [5:0]  pp343;
wire [5:0]  pp344;
wire [5:0]  pp345;
wire [5:0]  pp346;
wire [5:0]  pp347;
wire [5:0]  pp348;
wire [5:0]  pp349;
wire [5:0]  pp350;
wire [5:0]  pp351;
wire [5:0]  pp352;
wire [5:0]  pp353;
wire [5:0]  pp354;
wire [5:0]  pp355;
wire [5:0]  pp356;
wire [5:0]  pp357;
wire [5:0]  pp358;
wire [5:0]  pp359;
wire [5:0]  pp360;
wire [5:0]  pp361;
wire [5:0]  pp362;
wire [5:0]  pp363;
wire [5:0]  pp364;
wire [5:0]  pp365;
wire [5:0]  pp366;
wire [5:0]  pp367;
wire [5:0]  pp368;
wire [5:0]  pp369;
wire [5:0]  pp370;
wire [5:0]  pp371;
wire [5:0]  pp372;
wire [5:0]  pp373;
wire [5:0]  pp374;
wire [5:0]  pp375;
wire [5:0]  pp376;
wire [5:0]  pp377;
wire [5:0]  pp378;
wire [5:0]  pp379;
wire [5:0]  pp380;
wire [5:0]  pp381;
wire [5:0]  pp382;
wire [5:0]  pp383;
wire [5:0]  pp384;
wire [5:0]  pp385;
wire [5:0]  pp386;
wire [5:0]  pp387;
wire [5:0]  pp388;
wire [5:0]  pp389;
wire [5:0]  pp390;
wire [5:0]  pp391;
wire [5:0]  pp392;
wire [5:0]  pp393;
wire [5:0]  pp394;
wire [5:0]  pp395;
wire [5:0]  pp396;
wire [5:0]  pp397;
wire [5:0]  pp398;
wire [5:0]  pp399;
wire [5:0]  pp400;
wire [5:0]  pp401;
wire [5:0]  pp402;
wire [5:0]  pp403;
wire [5:0]  pp404;
wire [5:0]  pp405;
wire [5:0]  pp406;
wire [5:0]  pp407;
wire [5:0]  pp408;
wire [5:0]  pp409;
wire [5:0]  pp410;
wire [5:0]  pp411;
wire [5:0]  pp412;
wire [5:0]  pp413;
wire [5:0]  pp414;
wire [5:0]  pp415;
wire [5:0]  pp416;
wire [5:0]  pp417;
wire [5:0]  pp418;
wire [5:0]  pp419;
wire [5:0]  pp420;
wire [5:0]  pp421;
wire [5:0]  pp422;
wire [5:0]  pp423;
wire [5:0]  pp424;
wire [5:0]  pp425;
wire [5:0]  pp426;
wire [5:0]  pp427;
wire [5:0]  pp428;
wire [5:0]  pp429;
wire [5:0]  pp430;
wire [5:0]  pp431;
wire [5:0]  pp432;
wire [5:0]  pp433;
wire [5:0]  pp434;
wire [5:0]  pp435;
wire [5:0]  pp436;
wire [5:0]  pp437;
wire [5:0]  pp438;
wire [5:0]  pp439;
wire [5:0]  pp440;
wire [5:0]  pp441;
wire [5:0]  pp442;
wire [5:0]  pp443;
wire [5:0]  pp444;
wire [5:0]  pp445;
wire [5:0]  pp446;
wire [5:0]  pp447;
wire [5:0]  pp448;
wire [5:0]  pp449;
wire [5:0]  pp450;
wire [5:0]  pp451;
wire [5:0]  pp452;
wire [5:0]  pp453;
wire [5:0]  pp454;
wire [5:0]  pp455;
wire [5:0]  pp456;
wire [5:0]  pp457;
wire [5:0]  pp458;
wire [5:0]  pp459;
wire [5:0]  pp460;
wire [5:0]  pp461;
wire [5:0]  pp462;
wire [5:0]  pp463;
wire [5:0]  pp464;
wire [5:0]  pp465;
wire [5:0]  pp466;
wire [5:0]  pp467;
wire [5:0]  pp468;
wire [5:0]  pp469;
wire [5:0]  pp470;
wire [5:0]  pp471;
wire [5:0]  pp472;
wire [5:0]  pp473;
wire [5:0]  pp474;
wire [5:0]  pp475;
wire [5:0]  pp476;
wire [5:0]  pp477;
wire [5:0]  pp478;
wire [5:0]  pp479;
wire [5:0]  pp480;
wire [5:0]  pp481;
wire [5:0]  pp482;
wire [5:0]  pp483;
wire [5:0]  pp484;
wire [5:0]  pp485;
wire [5:0]  pp486;
wire [5:0]  pp487;
wire [5:0]  pp488;
wire [5:0]  pp489;
wire [5:0]  pp490;
wire [5:0]  pp491;
wire [5:0]  pp492;
wire [5:0]  pp493;
wire [5:0]  pp494;
wire [5:0]  pp495;
wire [5:0]  pp496;
wire [5:0]  pp497;
wire [5:0]  pp498;
wire [5:0]  pp499;
wire [5:0]  pp500;
wire [5:0]  pp501;
wire [5:0]  pp502;
wire [5:0]  pp503;
wire [5:0]  pp504;
wire [5:0]  pp505;
wire [5:0]  pp506;
wire [5:0]  pp507;
wire [5:0]  pp508;
wire [5:0]  pp509;
wire [5:0]  pp510;
wire [5:0]  pp511;

// partial products
level0_mult lvl0_mult0({in0[3:0], in1[1:0]}, pp0);
level0_mult lvl0_mult1({in0[7:4], in1[1:0]}, pp1);
level0_mult lvl0_mult2({in0[11:8], in1[1:0]}, pp2);
level0_mult lvl0_mult3({in0[15:12], in1[1:0]}, pp3);
level0_mult lvl0_mult4({in0[19:16], in1[1:0]}, pp4);
level0_mult lvl0_mult5({in0[23:20], in1[1:0]}, pp5);
level0_mult lvl0_mult6({in0[27:24], in1[1:0]}, pp6);
level0_mult lvl0_mult7({in0[31:28], in1[1:0]}, pp7);
level0_mult lvl0_mult8({in0[35:32], in1[1:0]}, pp8);
level0_mult lvl0_mult9({in0[39:36], in1[1:0]}, pp9);
level0_mult lvl0_mult10({in0[43:40], in1[1:0]}, pp10);
level0_mult lvl0_mult11({in0[47:44], in1[1:0]}, pp11);
level0_mult lvl0_mult12({in0[51:48], in1[1:0]}, pp12);
level0_mult lvl0_mult13({in0[55:52], in1[1:0]}, pp13);
level0_mult lvl0_mult14({in0[59:56], in1[1:0]}, pp14);
level0_mult lvl0_mult15({in0[63:60], in1[1:0]}, pp15);
level0_mult lvl0_mult16({in0[3:0], in1[3:2]}, pp16);
level0_mult lvl0_mult17({in0[7:4], in1[3:2]}, pp17);
level0_mult lvl0_mult18({in0[11:8], in1[3:2]}, pp18);
level0_mult lvl0_mult19({in0[15:12], in1[3:2]}, pp19);
level0_mult lvl0_mult20({in0[19:16], in1[3:2]}, pp20);
level0_mult lvl0_mult21({in0[23:20], in1[3:2]}, pp21);
level0_mult lvl0_mult22({in0[27:24], in1[3:2]}, pp22);
level0_mult lvl0_mult23({in0[31:28], in1[3:2]}, pp23);
level0_mult lvl0_mult24({in0[35:32], in1[3:2]}, pp24);
level0_mult lvl0_mult25({in0[39:36], in1[3:2]}, pp25);
level0_mult lvl0_mult26({in0[43:40], in1[3:2]}, pp26);
level0_mult lvl0_mult27({in0[47:44], in1[3:2]}, pp27);
level0_mult lvl0_mult28({in0[51:48], in1[3:2]}, pp28);
level0_mult lvl0_mult29({in0[55:52], in1[3:2]}, pp29);
level0_mult lvl0_mult30({in0[59:56], in1[3:2]}, pp30);
level0_mult lvl0_mult31({in0[63:60], in1[3:2]}, pp31);
level0_mult lvl0_mult32({in0[3:0], in1[5:4]}, pp32);
level0_mult lvl0_mult33({in0[7:4], in1[5:4]}, pp33);
level0_mult lvl0_mult34({in0[11:8], in1[5:4]}, pp34);
level0_mult lvl0_mult35({in0[15:12], in1[5:4]}, pp35);
level0_mult lvl0_mult36({in0[19:16], in1[5:4]}, pp36);
level0_mult lvl0_mult37({in0[23:20], in1[5:4]}, pp37);
level0_mult lvl0_mult38({in0[27:24], in1[5:4]}, pp38);
level0_mult lvl0_mult39({in0[31:28], in1[5:4]}, pp39);
level0_mult lvl0_mult40({in0[35:32], in1[5:4]}, pp40);
level0_mult lvl0_mult41({in0[39:36], in1[5:4]}, pp41);
level0_mult lvl0_mult42({in0[43:40], in1[5:4]}, pp42);
level0_mult lvl0_mult43({in0[47:44], in1[5:4]}, pp43);
level0_mult lvl0_mult44({in0[51:48], in1[5:4]}, pp44);
level0_mult lvl0_mult45({in0[55:52], in1[5:4]}, pp45);
level0_mult lvl0_mult46({in0[59:56], in1[5:4]}, pp46);
level0_mult lvl0_mult47({in0[63:60], in1[5:4]}, pp47);
level0_mult lvl0_mult48({in0[3:0], in1[7:6]}, pp48);
level0_mult lvl0_mult49({in0[7:4], in1[7:6]}, pp49);
level0_mult lvl0_mult50({in0[11:8], in1[7:6]}, pp50);
level0_mult lvl0_mult51({in0[15:12], in1[7:6]}, pp51);
level0_mult lvl0_mult52({in0[19:16], in1[7:6]}, pp52);
level0_mult lvl0_mult53({in0[23:20], in1[7:6]}, pp53);
level0_mult lvl0_mult54({in0[27:24], in1[7:6]}, pp54);
level0_mult lvl0_mult55({in0[31:28], in1[7:6]}, pp55);
level0_mult lvl0_mult56({in0[35:32], in1[7:6]}, pp56);
level0_mult lvl0_mult57({in0[39:36], in1[7:6]}, pp57);
level0_mult lvl0_mult58({in0[43:40], in1[7:6]}, pp58);
level0_mult lvl0_mult59({in0[47:44], in1[7:6]}, pp59);
level0_mult lvl0_mult60({in0[51:48], in1[7:6]}, pp60);
level0_mult lvl0_mult61({in0[55:52], in1[7:6]}, pp61);
level0_mult lvl0_mult62({in0[59:56], in1[7:6]}, pp62);
level0_mult lvl0_mult63({in0[63:60], in1[7:6]}, pp63);
level0_mult lvl0_mult64({in0[3:0], in1[9:8]}, pp64);
level0_mult lvl0_mult65({in0[7:4], in1[9:8]}, pp65);
level0_mult lvl0_mult66({in0[11:8], in1[9:8]}, pp66);
level0_mult lvl0_mult67({in0[15:12], in1[9:8]}, pp67);
level0_mult lvl0_mult68({in0[19:16], in1[9:8]}, pp68);
level0_mult lvl0_mult69({in0[23:20], in1[9:8]}, pp69);
level0_mult lvl0_mult70({in0[27:24], in1[9:8]}, pp70);
level0_mult lvl0_mult71({in0[31:28], in1[9:8]}, pp71);
level0_mult lvl0_mult72({in0[35:32], in1[9:8]}, pp72);
level0_mult lvl0_mult73({in0[39:36], in1[9:8]}, pp73);
level0_mult lvl0_mult74({in0[43:40], in1[9:8]}, pp74);
level0_mult lvl0_mult75({in0[47:44], in1[9:8]}, pp75);
level0_mult lvl0_mult76({in0[51:48], in1[9:8]}, pp76);
level0_mult lvl0_mult77({in0[55:52], in1[9:8]}, pp77);
level0_mult lvl0_mult78({in0[59:56], in1[9:8]}, pp78);
level0_mult lvl0_mult79({in0[63:60], in1[9:8]}, pp79);
level0_mult lvl0_mult80({in0[3:0], in1[11:10]}, pp80);
level0_mult lvl0_mult81({in0[7:4], in1[11:10]}, pp81);
level0_mult lvl0_mult82({in0[11:8], in1[11:10]}, pp82);
level0_mult lvl0_mult83({in0[15:12], in1[11:10]}, pp83);
level0_mult lvl0_mult84({in0[19:16], in1[11:10]}, pp84);
level0_mult lvl0_mult85({in0[23:20], in1[11:10]}, pp85);
level0_mult lvl0_mult86({in0[27:24], in1[11:10]}, pp86);
level0_mult lvl0_mult87({in0[31:28], in1[11:10]}, pp87);
level0_mult lvl0_mult88({in0[35:32], in1[11:10]}, pp88);
level0_mult lvl0_mult89({in0[39:36], in1[11:10]}, pp89);
level0_mult lvl0_mult90({in0[43:40], in1[11:10]}, pp90);
level0_mult lvl0_mult91({in0[47:44], in1[11:10]}, pp91);
level0_mult lvl0_mult92({in0[51:48], in1[11:10]}, pp92);
level0_mult lvl0_mult93({in0[55:52], in1[11:10]}, pp93);
level0_mult lvl0_mult94({in0[59:56], in1[11:10]}, pp94);
level0_mult lvl0_mult95({in0[63:60], in1[11:10]}, pp95);
level0_mult lvl0_mult96({in0[3:0], in1[13:12]}, pp96);
level0_mult lvl0_mult97({in0[7:4], in1[13:12]}, pp97);
level0_mult lvl0_mult98({in0[11:8], in1[13:12]}, pp98);
level0_mult lvl0_mult99({in0[15:12], in1[13:12]}, pp99);
level0_mult lvl0_mult100({in0[19:16], in1[13:12]}, pp100);
level0_mult lvl0_mult101({in0[23:20], in1[13:12]}, pp101);
level0_mult lvl0_mult102({in0[27:24], in1[13:12]}, pp102);
level0_mult lvl0_mult103({in0[31:28], in1[13:12]}, pp103);
level0_mult lvl0_mult104({in0[35:32], in1[13:12]}, pp104);
level0_mult lvl0_mult105({in0[39:36], in1[13:12]}, pp105);
level0_mult lvl0_mult106({in0[43:40], in1[13:12]}, pp106);
level0_mult lvl0_mult107({in0[47:44], in1[13:12]}, pp107);
level0_mult lvl0_mult108({in0[51:48], in1[13:12]}, pp108);
level0_mult lvl0_mult109({in0[55:52], in1[13:12]}, pp109);
level0_mult lvl0_mult110({in0[59:56], in1[13:12]}, pp110);
level0_mult lvl0_mult111({in0[63:60], in1[13:12]}, pp111);
level0_mult lvl0_mult112({in0[3:0], in1[15:14]}, pp112);
level0_mult lvl0_mult113({in0[7:4], in1[15:14]}, pp113);
level0_mult lvl0_mult114({in0[11:8], in1[15:14]}, pp114);
level0_mult lvl0_mult115({in0[15:12], in1[15:14]}, pp115);
level0_mult lvl0_mult116({in0[19:16], in1[15:14]}, pp116);
level0_mult lvl0_mult117({in0[23:20], in1[15:14]}, pp117);
level0_mult lvl0_mult118({in0[27:24], in1[15:14]}, pp118);
level0_mult lvl0_mult119({in0[31:28], in1[15:14]}, pp119);
level0_mult lvl0_mult120({in0[35:32], in1[15:14]}, pp120);
level0_mult lvl0_mult121({in0[39:36], in1[15:14]}, pp121);
level0_mult lvl0_mult122({in0[43:40], in1[15:14]}, pp122);
level0_mult lvl0_mult123({in0[47:44], in1[15:14]}, pp123);
level0_mult lvl0_mult124({in0[51:48], in1[15:14]}, pp124);
level0_mult lvl0_mult125({in0[55:52], in1[15:14]}, pp125);
level0_mult lvl0_mult126({in0[59:56], in1[15:14]}, pp126);
level0_mult lvl0_mult127({in0[63:60], in1[15:14]}, pp127);
level0_mult lvl0_mult128({in0[3:0], in1[17:16]}, pp128);
level0_mult lvl0_mult129({in0[7:4], in1[17:16]}, pp129);
level0_mult lvl0_mult130({in0[11:8], in1[17:16]}, pp130);
level0_mult lvl0_mult131({in0[15:12], in1[17:16]}, pp131);
level0_mult lvl0_mult132({in0[19:16], in1[17:16]}, pp132);
level0_mult lvl0_mult133({in0[23:20], in1[17:16]}, pp133);
level0_mult lvl0_mult134({in0[27:24], in1[17:16]}, pp134);
level0_mult lvl0_mult135({in0[31:28], in1[17:16]}, pp135);
level0_mult lvl0_mult136({in0[35:32], in1[17:16]}, pp136);
level0_mult lvl0_mult137({in0[39:36], in1[17:16]}, pp137);
level0_mult lvl0_mult138({in0[43:40], in1[17:16]}, pp138);
level0_mult lvl0_mult139({in0[47:44], in1[17:16]}, pp139);
level0_mult lvl0_mult140({in0[51:48], in1[17:16]}, pp140);
level0_mult lvl0_mult141({in0[55:52], in1[17:16]}, pp141);
level0_mult lvl0_mult142({in0[59:56], in1[17:16]}, pp142);
level0_mult lvl0_mult143({in0[63:60], in1[17:16]}, pp143);
level0_mult lvl0_mult144({in0[3:0], in1[19:18]}, pp144);
level0_mult lvl0_mult145({in0[7:4], in1[19:18]}, pp145);
level0_mult lvl0_mult146({in0[11:8], in1[19:18]}, pp146);
level0_mult lvl0_mult147({in0[15:12], in1[19:18]}, pp147);
level0_mult lvl0_mult148({in0[19:16], in1[19:18]}, pp148);
level0_mult lvl0_mult149({in0[23:20], in1[19:18]}, pp149);
level0_mult lvl0_mult150({in0[27:24], in1[19:18]}, pp150);
level0_mult lvl0_mult151({in0[31:28], in1[19:18]}, pp151);
level0_mult lvl0_mult152({in0[35:32], in1[19:18]}, pp152);
level0_mult lvl0_mult153({in0[39:36], in1[19:18]}, pp153);
level0_mult lvl0_mult154({in0[43:40], in1[19:18]}, pp154);
level0_mult lvl0_mult155({in0[47:44], in1[19:18]}, pp155);
level0_mult lvl0_mult156({in0[51:48], in1[19:18]}, pp156);
level0_mult lvl0_mult157({in0[55:52], in1[19:18]}, pp157);
level0_mult lvl0_mult158({in0[59:56], in1[19:18]}, pp158);
level0_mult lvl0_mult159({in0[63:60], in1[19:18]}, pp159);
level0_mult lvl0_mult160({in0[3:0], in1[21:20]}, pp160);
level0_mult lvl0_mult161({in0[7:4], in1[21:20]}, pp161);
level0_mult lvl0_mult162({in0[11:8], in1[21:20]}, pp162);
level0_mult lvl0_mult163({in0[15:12], in1[21:20]}, pp163);
level0_mult lvl0_mult164({in0[19:16], in1[21:20]}, pp164);
level0_mult lvl0_mult165({in0[23:20], in1[21:20]}, pp165);
level0_mult lvl0_mult166({in0[27:24], in1[21:20]}, pp166);
level0_mult lvl0_mult167({in0[31:28], in1[21:20]}, pp167);
level0_mult lvl0_mult168({in0[35:32], in1[21:20]}, pp168);
level0_mult lvl0_mult169({in0[39:36], in1[21:20]}, pp169);
level0_mult lvl0_mult170({in0[43:40], in1[21:20]}, pp170);
level0_mult lvl0_mult171({in0[47:44], in1[21:20]}, pp171);
level0_mult lvl0_mult172({in0[51:48], in1[21:20]}, pp172);
level0_mult lvl0_mult173({in0[55:52], in1[21:20]}, pp173);
level0_mult lvl0_mult174({in0[59:56], in1[21:20]}, pp174);
level0_mult lvl0_mult175({in0[63:60], in1[21:20]}, pp175);
level0_mult lvl0_mult176({in0[3:0], in1[23:22]}, pp176);
level0_mult lvl0_mult177({in0[7:4], in1[23:22]}, pp177);
level0_mult lvl0_mult178({in0[11:8], in1[23:22]}, pp178);
level0_mult lvl0_mult179({in0[15:12], in1[23:22]}, pp179);
level0_mult lvl0_mult180({in0[19:16], in1[23:22]}, pp180);
level0_mult lvl0_mult181({in0[23:20], in1[23:22]}, pp181);
level0_mult lvl0_mult182({in0[27:24], in1[23:22]}, pp182);
level0_mult lvl0_mult183({in0[31:28], in1[23:22]}, pp183);
level0_mult lvl0_mult184({in0[35:32], in1[23:22]}, pp184);
level0_mult lvl0_mult185({in0[39:36], in1[23:22]}, pp185);
level0_mult lvl0_mult186({in0[43:40], in1[23:22]}, pp186);
level0_mult lvl0_mult187({in0[47:44], in1[23:22]}, pp187);
level0_mult lvl0_mult188({in0[51:48], in1[23:22]}, pp188);
level0_mult lvl0_mult189({in0[55:52], in1[23:22]}, pp189);
level0_mult lvl0_mult190({in0[59:56], in1[23:22]}, pp190);
level0_mult lvl0_mult191({in0[63:60], in1[23:22]}, pp191);
level0_mult lvl0_mult192({in0[3:0], in1[25:24]}, pp192);
level0_mult lvl0_mult193({in0[7:4], in1[25:24]}, pp193);
level0_mult lvl0_mult194({in0[11:8], in1[25:24]}, pp194);
level0_mult lvl0_mult195({in0[15:12], in1[25:24]}, pp195);
level0_mult lvl0_mult196({in0[19:16], in1[25:24]}, pp196);
level0_mult lvl0_mult197({in0[23:20], in1[25:24]}, pp197);
level0_mult lvl0_mult198({in0[27:24], in1[25:24]}, pp198);
level0_mult lvl0_mult199({in0[31:28], in1[25:24]}, pp199);
level0_mult lvl0_mult200({in0[35:32], in1[25:24]}, pp200);
level0_mult lvl0_mult201({in0[39:36], in1[25:24]}, pp201);
level0_mult lvl0_mult202({in0[43:40], in1[25:24]}, pp202);
level0_mult lvl0_mult203({in0[47:44], in1[25:24]}, pp203);
level0_mult lvl0_mult204({in0[51:48], in1[25:24]}, pp204);
level0_mult lvl0_mult205({in0[55:52], in1[25:24]}, pp205);
level0_mult lvl0_mult206({in0[59:56], in1[25:24]}, pp206);
level0_mult lvl0_mult207({in0[63:60], in1[25:24]}, pp207);
level0_mult lvl0_mult208({in0[3:0], in1[27:26]}, pp208);
level0_mult lvl0_mult209({in0[7:4], in1[27:26]}, pp209);
level0_mult lvl0_mult210({in0[11:8], in1[27:26]}, pp210);
level0_mult lvl0_mult211({in0[15:12], in1[27:26]}, pp211);
level0_mult lvl0_mult212({in0[19:16], in1[27:26]}, pp212);
level0_mult lvl0_mult213({in0[23:20], in1[27:26]}, pp213);
level0_mult lvl0_mult214({in0[27:24], in1[27:26]}, pp214);
level0_mult lvl0_mult215({in0[31:28], in1[27:26]}, pp215);
level0_mult lvl0_mult216({in0[35:32], in1[27:26]}, pp216);
level0_mult lvl0_mult217({in0[39:36], in1[27:26]}, pp217);
level0_mult lvl0_mult218({in0[43:40], in1[27:26]}, pp218);
level0_mult lvl0_mult219({in0[47:44], in1[27:26]}, pp219);
level0_mult lvl0_mult220({in0[51:48], in1[27:26]}, pp220);
level0_mult lvl0_mult221({in0[55:52], in1[27:26]}, pp221);
level0_mult lvl0_mult222({in0[59:56], in1[27:26]}, pp222);
level0_mult lvl0_mult223({in0[63:60], in1[27:26]}, pp223);
level0_mult lvl0_mult224({in0[3:0], in1[29:28]}, pp224);
level0_mult lvl0_mult225({in0[7:4], in1[29:28]}, pp225);
level0_mult lvl0_mult226({in0[11:8], in1[29:28]}, pp226);
level0_mult lvl0_mult227({in0[15:12], in1[29:28]}, pp227);
level0_mult lvl0_mult228({in0[19:16], in1[29:28]}, pp228);
level0_mult lvl0_mult229({in0[23:20], in1[29:28]}, pp229);
level0_mult lvl0_mult230({in0[27:24], in1[29:28]}, pp230);
level0_mult lvl0_mult231({in0[31:28], in1[29:28]}, pp231);
level0_mult lvl0_mult232({in0[35:32], in1[29:28]}, pp232);
level0_mult lvl0_mult233({in0[39:36], in1[29:28]}, pp233);
level0_mult lvl0_mult234({in0[43:40], in1[29:28]}, pp234);
level0_mult lvl0_mult235({in0[47:44], in1[29:28]}, pp235);
level0_mult lvl0_mult236({in0[51:48], in1[29:28]}, pp236);
level0_mult lvl0_mult237({in0[55:52], in1[29:28]}, pp237);
level0_mult lvl0_mult238({in0[59:56], in1[29:28]}, pp238);
level0_mult lvl0_mult239({in0[63:60], in1[29:28]}, pp239);
level0_mult lvl0_mult240({in0[3:0], in1[31:30]}, pp240);
level0_mult lvl0_mult241({in0[7:4], in1[31:30]}, pp241);
level0_mult lvl0_mult242({in0[11:8], in1[31:30]}, pp242);
level0_mult lvl0_mult243({in0[15:12], in1[31:30]}, pp243);
level0_mult lvl0_mult244({in0[19:16], in1[31:30]}, pp244);
level0_mult lvl0_mult245({in0[23:20], in1[31:30]}, pp245);
level0_mult lvl0_mult246({in0[27:24], in1[31:30]}, pp246);
level0_mult lvl0_mult247({in0[31:28], in1[31:30]}, pp247);
level0_mult lvl0_mult248({in0[35:32], in1[31:30]}, pp248);
level0_mult lvl0_mult249({in0[39:36], in1[31:30]}, pp249);
level0_mult lvl0_mult250({in0[43:40], in1[31:30]}, pp250);
level0_mult lvl0_mult251({in0[47:44], in1[31:30]}, pp251);
level0_mult lvl0_mult252({in0[51:48], in1[31:30]}, pp252);
level0_mult lvl0_mult253({in0[55:52], in1[31:30]}, pp253);
level0_mult lvl0_mult254({in0[59:56], in1[31:30]}, pp254);
level0_mult lvl0_mult255({in0[63:60], in1[31:30]}, pp255);
level0_mult lvl0_mult256({in0[3:0], in1[33:32]}, pp256);
level0_mult lvl0_mult257({in0[7:4], in1[33:32]}, pp257);
level0_mult lvl0_mult258({in0[11:8], in1[33:32]}, pp258);
level0_mult lvl0_mult259({in0[15:12], in1[33:32]}, pp259);
level0_mult lvl0_mult260({in0[19:16], in1[33:32]}, pp260);
level0_mult lvl0_mult261({in0[23:20], in1[33:32]}, pp261);
level0_mult lvl0_mult262({in0[27:24], in1[33:32]}, pp262);
level0_mult lvl0_mult263({in0[31:28], in1[33:32]}, pp263);
level0_mult lvl0_mult264({in0[35:32], in1[33:32]}, pp264);
level0_mult lvl0_mult265({in0[39:36], in1[33:32]}, pp265);
level0_mult lvl0_mult266({in0[43:40], in1[33:32]}, pp266);
level0_mult lvl0_mult267({in0[47:44], in1[33:32]}, pp267);
level0_mult lvl0_mult268({in0[51:48], in1[33:32]}, pp268);
level0_mult lvl0_mult269({in0[55:52], in1[33:32]}, pp269);
level0_mult lvl0_mult270({in0[59:56], in1[33:32]}, pp270);
level0_mult lvl0_mult271({in0[63:60], in1[33:32]}, pp271);
level0_mult lvl0_mult272({in0[3:0], in1[35:34]}, pp272);
level0_mult lvl0_mult273({in0[7:4], in1[35:34]}, pp273);
level0_mult lvl0_mult274({in0[11:8], in1[35:34]}, pp274);
level0_mult lvl0_mult275({in0[15:12], in1[35:34]}, pp275);
level0_mult lvl0_mult276({in0[19:16], in1[35:34]}, pp276);
level0_mult lvl0_mult277({in0[23:20], in1[35:34]}, pp277);
level0_mult lvl0_mult278({in0[27:24], in1[35:34]}, pp278);
level0_mult lvl0_mult279({in0[31:28], in1[35:34]}, pp279);
level0_mult lvl0_mult280({in0[35:32], in1[35:34]}, pp280);
level0_mult lvl0_mult281({in0[39:36], in1[35:34]}, pp281);
level0_mult lvl0_mult282({in0[43:40], in1[35:34]}, pp282);
level0_mult lvl0_mult283({in0[47:44], in1[35:34]}, pp283);
level0_mult lvl0_mult284({in0[51:48], in1[35:34]}, pp284);
level0_mult lvl0_mult285({in0[55:52], in1[35:34]}, pp285);
level0_mult lvl0_mult286({in0[59:56], in1[35:34]}, pp286);
level0_mult lvl0_mult287({in0[63:60], in1[35:34]}, pp287);
level0_mult lvl0_mult288({in0[3:0], in1[37:36]}, pp288);
level0_mult lvl0_mult289({in0[7:4], in1[37:36]}, pp289);
level0_mult lvl0_mult290({in0[11:8], in1[37:36]}, pp290);
level0_mult lvl0_mult291({in0[15:12], in1[37:36]}, pp291);
level0_mult lvl0_mult292({in0[19:16], in1[37:36]}, pp292);
level0_mult lvl0_mult293({in0[23:20], in1[37:36]}, pp293);
level0_mult lvl0_mult294({in0[27:24], in1[37:36]}, pp294);
level0_mult lvl0_mult295({in0[31:28], in1[37:36]}, pp295);
level0_mult lvl0_mult296({in0[35:32], in1[37:36]}, pp296);
level0_mult lvl0_mult297({in0[39:36], in1[37:36]}, pp297);
level0_mult lvl0_mult298({in0[43:40], in1[37:36]}, pp298);
level0_mult lvl0_mult299({in0[47:44], in1[37:36]}, pp299);
level0_mult lvl0_mult300({in0[51:48], in1[37:36]}, pp300);
level0_mult lvl0_mult301({in0[55:52], in1[37:36]}, pp301);
level0_mult lvl0_mult302({in0[59:56], in1[37:36]}, pp302);
level0_mult lvl0_mult303({in0[63:60], in1[37:36]}, pp303);
level0_mult lvl0_mult304({in0[3:0], in1[39:38]}, pp304);
level0_mult lvl0_mult305({in0[7:4], in1[39:38]}, pp305);
level0_mult lvl0_mult306({in0[11:8], in1[39:38]}, pp306);
level0_mult lvl0_mult307({in0[15:12], in1[39:38]}, pp307);
level0_mult lvl0_mult308({in0[19:16], in1[39:38]}, pp308);
level0_mult lvl0_mult309({in0[23:20], in1[39:38]}, pp309);
level0_mult lvl0_mult310({in0[27:24], in1[39:38]}, pp310);
level0_mult lvl0_mult311({in0[31:28], in1[39:38]}, pp311);
level0_mult lvl0_mult312({in0[35:32], in1[39:38]}, pp312);
level0_mult lvl0_mult313({in0[39:36], in1[39:38]}, pp313);
level0_mult lvl0_mult314({in0[43:40], in1[39:38]}, pp314);
level0_mult lvl0_mult315({in0[47:44], in1[39:38]}, pp315);
level0_mult lvl0_mult316({in0[51:48], in1[39:38]}, pp316);
level0_mult lvl0_mult317({in0[55:52], in1[39:38]}, pp317);
level0_mult lvl0_mult318({in0[59:56], in1[39:38]}, pp318);
level0_mult lvl0_mult319({in0[63:60], in1[39:38]}, pp319);
level0_mult lvl0_mult320({in0[3:0], in1[41:40]}, pp320);
level0_mult lvl0_mult321({in0[7:4], in1[41:40]}, pp321);
level0_mult lvl0_mult322({in0[11:8], in1[41:40]}, pp322);
level0_mult lvl0_mult323({in0[15:12], in1[41:40]}, pp323);
level0_mult lvl0_mult324({in0[19:16], in1[41:40]}, pp324);
level0_mult lvl0_mult325({in0[23:20], in1[41:40]}, pp325);
level0_mult lvl0_mult326({in0[27:24], in1[41:40]}, pp326);
level0_mult lvl0_mult327({in0[31:28], in1[41:40]}, pp327);
level0_mult lvl0_mult328({in0[35:32], in1[41:40]}, pp328);
level0_mult lvl0_mult329({in0[39:36], in1[41:40]}, pp329);
level0_mult lvl0_mult330({in0[43:40], in1[41:40]}, pp330);
level0_mult lvl0_mult331({in0[47:44], in1[41:40]}, pp331);
level0_mult lvl0_mult332({in0[51:48], in1[41:40]}, pp332);
level0_mult lvl0_mult333({in0[55:52], in1[41:40]}, pp333);
level0_mult lvl0_mult334({in0[59:56], in1[41:40]}, pp334);
level0_mult lvl0_mult335({in0[63:60], in1[41:40]}, pp335);
level0_mult lvl0_mult336({in0[3:0], in1[43:42]}, pp336);
level0_mult lvl0_mult337({in0[7:4], in1[43:42]}, pp337);
level0_mult lvl0_mult338({in0[11:8], in1[43:42]}, pp338);
level0_mult lvl0_mult339({in0[15:12], in1[43:42]}, pp339);
level0_mult lvl0_mult340({in0[19:16], in1[43:42]}, pp340);
level0_mult lvl0_mult341({in0[23:20], in1[43:42]}, pp341);
level0_mult lvl0_mult342({in0[27:24], in1[43:42]}, pp342);
level0_mult lvl0_mult343({in0[31:28], in1[43:42]}, pp343);
level0_mult lvl0_mult344({in0[35:32], in1[43:42]}, pp344);
level0_mult lvl0_mult345({in0[39:36], in1[43:42]}, pp345);
level0_mult lvl0_mult346({in0[43:40], in1[43:42]}, pp346);
level0_mult lvl0_mult347({in0[47:44], in1[43:42]}, pp347);
level0_mult lvl0_mult348({in0[51:48], in1[43:42]}, pp348);
level0_mult lvl0_mult349({in0[55:52], in1[43:42]}, pp349);
level0_mult lvl0_mult350({in0[59:56], in1[43:42]}, pp350);
level0_mult lvl0_mult351({in0[63:60], in1[43:42]}, pp351);
level0_mult lvl0_mult352({in0[3:0], in1[45:44]}, pp352);
level0_mult lvl0_mult353({in0[7:4], in1[45:44]}, pp353);
level0_mult lvl0_mult354({in0[11:8], in1[45:44]}, pp354);
level0_mult lvl0_mult355({in0[15:12], in1[45:44]}, pp355);
level0_mult lvl0_mult356({in0[19:16], in1[45:44]}, pp356);
level0_mult lvl0_mult357({in0[23:20], in1[45:44]}, pp357);
level0_mult lvl0_mult358({in0[27:24], in1[45:44]}, pp358);
level0_mult lvl0_mult359({in0[31:28], in1[45:44]}, pp359);
level0_mult lvl0_mult360({in0[35:32], in1[45:44]}, pp360);
level0_mult lvl0_mult361({in0[39:36], in1[45:44]}, pp361);
level0_mult lvl0_mult362({in0[43:40], in1[45:44]}, pp362);
level0_mult lvl0_mult363({in0[47:44], in1[45:44]}, pp363);
level0_mult lvl0_mult364({in0[51:48], in1[45:44]}, pp364);
level0_mult lvl0_mult365({in0[55:52], in1[45:44]}, pp365);
level0_mult lvl0_mult366({in0[59:56], in1[45:44]}, pp366);
level0_mult lvl0_mult367({in0[63:60], in1[45:44]}, pp367);
level0_mult lvl0_mult368({in0[3:0], in1[47:46]}, pp368);
level0_mult lvl0_mult369({in0[7:4], in1[47:46]}, pp369);
level0_mult lvl0_mult370({in0[11:8], in1[47:46]}, pp370);
level0_mult lvl0_mult371({in0[15:12], in1[47:46]}, pp371);
level0_mult lvl0_mult372({in0[19:16], in1[47:46]}, pp372);
level0_mult lvl0_mult373({in0[23:20], in1[47:46]}, pp373);
level0_mult lvl0_mult374({in0[27:24], in1[47:46]}, pp374);
level0_mult lvl0_mult375({in0[31:28], in1[47:46]}, pp375);
level0_mult lvl0_mult376({in0[35:32], in1[47:46]}, pp376);
level0_mult lvl0_mult377({in0[39:36], in1[47:46]}, pp377);
level0_mult lvl0_mult378({in0[43:40], in1[47:46]}, pp378);
level0_mult lvl0_mult379({in0[47:44], in1[47:46]}, pp379);
level0_mult lvl0_mult380({in0[51:48], in1[47:46]}, pp380);
level0_mult lvl0_mult381({in0[55:52], in1[47:46]}, pp381);
level0_mult lvl0_mult382({in0[59:56], in1[47:46]}, pp382);
level0_mult lvl0_mult383({in0[63:60], in1[47:46]}, pp383);
level0_mult lvl0_mult384({in0[3:0], in1[49:48]}, pp384);
level0_mult lvl0_mult385({in0[7:4], in1[49:48]}, pp385);
level0_mult lvl0_mult386({in0[11:8], in1[49:48]}, pp386);
level0_mult lvl0_mult387({in0[15:12], in1[49:48]}, pp387);
level0_mult lvl0_mult388({in0[19:16], in1[49:48]}, pp388);
level0_mult lvl0_mult389({in0[23:20], in1[49:48]}, pp389);
level0_mult lvl0_mult390({in0[27:24], in1[49:48]}, pp390);
level0_mult lvl0_mult391({in0[31:28], in1[49:48]}, pp391);
level0_mult lvl0_mult392({in0[35:32], in1[49:48]}, pp392);
level0_mult lvl0_mult393({in0[39:36], in1[49:48]}, pp393);
level0_mult lvl0_mult394({in0[43:40], in1[49:48]}, pp394);
level0_mult lvl0_mult395({in0[47:44], in1[49:48]}, pp395);
level0_mult lvl0_mult396({in0[51:48], in1[49:48]}, pp396);
level0_mult lvl0_mult397({in0[55:52], in1[49:48]}, pp397);
level0_mult lvl0_mult398({in0[59:56], in1[49:48]}, pp398);
level0_mult lvl0_mult399({in0[63:60], in1[49:48]}, pp399);
level0_mult lvl0_mult400({in0[3:0], in1[51:50]}, pp400);
level0_mult lvl0_mult401({in0[7:4], in1[51:50]}, pp401);
level0_mult lvl0_mult402({in0[11:8], in1[51:50]}, pp402);
level0_mult lvl0_mult403({in0[15:12], in1[51:50]}, pp403);
level0_mult lvl0_mult404({in0[19:16], in1[51:50]}, pp404);
level0_mult lvl0_mult405({in0[23:20], in1[51:50]}, pp405);
level0_mult lvl0_mult406({in0[27:24], in1[51:50]}, pp406);
level0_mult lvl0_mult407({in0[31:28], in1[51:50]}, pp407);
level0_mult lvl0_mult408({in0[35:32], in1[51:50]}, pp408);
level0_mult lvl0_mult409({in0[39:36], in1[51:50]}, pp409);
level0_mult lvl0_mult410({in0[43:40], in1[51:50]}, pp410);
level0_mult lvl0_mult411({in0[47:44], in1[51:50]}, pp411);
level0_mult lvl0_mult412({in0[51:48], in1[51:50]}, pp412);
level0_mult lvl0_mult413({in0[55:52], in1[51:50]}, pp413);
level0_mult lvl0_mult414({in0[59:56], in1[51:50]}, pp414);
level0_mult lvl0_mult415({in0[63:60], in1[51:50]}, pp415);
level0_mult lvl0_mult416({in0[3:0], in1[53:52]}, pp416);
level0_mult lvl0_mult417({in0[7:4], in1[53:52]}, pp417);
level0_mult lvl0_mult418({in0[11:8], in1[53:52]}, pp418);
level0_mult lvl0_mult419({in0[15:12], in1[53:52]}, pp419);
level0_mult lvl0_mult420({in0[19:16], in1[53:52]}, pp420);
level0_mult lvl0_mult421({in0[23:20], in1[53:52]}, pp421);
level0_mult lvl0_mult422({in0[27:24], in1[53:52]}, pp422);
level0_mult lvl0_mult423({in0[31:28], in1[53:52]}, pp423);
level0_mult lvl0_mult424({in0[35:32], in1[53:52]}, pp424);
level0_mult lvl0_mult425({in0[39:36], in1[53:52]}, pp425);
level0_mult lvl0_mult426({in0[43:40], in1[53:52]}, pp426);
level0_mult lvl0_mult427({in0[47:44], in1[53:52]}, pp427);
level0_mult lvl0_mult428({in0[51:48], in1[53:52]}, pp428);
level0_mult lvl0_mult429({in0[55:52], in1[53:52]}, pp429);
level0_mult lvl0_mult430({in0[59:56], in1[53:52]}, pp430);
level0_mult lvl0_mult431({in0[63:60], in1[53:52]}, pp431);
level0_mult lvl0_mult432({in0[3:0], in1[55:54]}, pp432);
level0_mult lvl0_mult433({in0[7:4], in1[55:54]}, pp433);
level0_mult lvl0_mult434({in0[11:8], in1[55:54]}, pp434);
level0_mult lvl0_mult435({in0[15:12], in1[55:54]}, pp435);
level0_mult lvl0_mult436({in0[19:16], in1[55:54]}, pp436);
level0_mult lvl0_mult437({in0[23:20], in1[55:54]}, pp437);
level0_mult lvl0_mult438({in0[27:24], in1[55:54]}, pp438);
level0_mult lvl0_mult439({in0[31:28], in1[55:54]}, pp439);
level0_mult lvl0_mult440({in0[35:32], in1[55:54]}, pp440);
level0_mult lvl0_mult441({in0[39:36], in1[55:54]}, pp441);
level0_mult lvl0_mult442({in0[43:40], in1[55:54]}, pp442);
level0_mult lvl0_mult443({in0[47:44], in1[55:54]}, pp443);
level0_mult lvl0_mult444({in0[51:48], in1[55:54]}, pp444);
level0_mult lvl0_mult445({in0[55:52], in1[55:54]}, pp445);
level0_mult lvl0_mult446({in0[59:56], in1[55:54]}, pp446);
level0_mult lvl0_mult447({in0[63:60], in1[55:54]}, pp447);
level0_mult lvl0_mult448({in0[3:0], in1[57:56]}, pp448);
level0_mult lvl0_mult449({in0[7:4], in1[57:56]}, pp449);
level0_mult lvl0_mult450({in0[11:8], in1[57:56]}, pp450);
level0_mult lvl0_mult451({in0[15:12], in1[57:56]}, pp451);
level0_mult lvl0_mult452({in0[19:16], in1[57:56]}, pp452);
level0_mult lvl0_mult453({in0[23:20], in1[57:56]}, pp453);
level0_mult lvl0_mult454({in0[27:24], in1[57:56]}, pp454);
level0_mult lvl0_mult455({in0[31:28], in1[57:56]}, pp455);
level0_mult lvl0_mult456({in0[35:32], in1[57:56]}, pp456);
level0_mult lvl0_mult457({in0[39:36], in1[57:56]}, pp457);
level0_mult lvl0_mult458({in0[43:40], in1[57:56]}, pp458);
level0_mult lvl0_mult459({in0[47:44], in1[57:56]}, pp459);
level0_mult lvl0_mult460({in0[51:48], in1[57:56]}, pp460);
level0_mult lvl0_mult461({in0[55:52], in1[57:56]}, pp461);
level0_mult lvl0_mult462({in0[59:56], in1[57:56]}, pp462);
level0_mult lvl0_mult463({in0[63:60], in1[57:56]}, pp463);
level0_mult lvl0_mult464({in0[3:0], in1[59:58]}, pp464);
level0_mult lvl0_mult465({in0[7:4], in1[59:58]}, pp465);
level0_mult lvl0_mult466({in0[11:8], in1[59:58]}, pp466);
level0_mult lvl0_mult467({in0[15:12], in1[59:58]}, pp467);
level0_mult lvl0_mult468({in0[19:16], in1[59:58]}, pp468);
level0_mult lvl0_mult469({in0[23:20], in1[59:58]}, pp469);
level0_mult lvl0_mult470({in0[27:24], in1[59:58]}, pp470);
level0_mult lvl0_mult471({in0[31:28], in1[59:58]}, pp471);
level0_mult lvl0_mult472({in0[35:32], in1[59:58]}, pp472);
level0_mult lvl0_mult473({in0[39:36], in1[59:58]}, pp473);
level0_mult lvl0_mult474({in0[43:40], in1[59:58]}, pp474);
level0_mult lvl0_mult475({in0[47:44], in1[59:58]}, pp475);
level0_mult lvl0_mult476({in0[51:48], in1[59:58]}, pp476);
level0_mult lvl0_mult477({in0[55:52], in1[59:58]}, pp477);
level0_mult lvl0_mult478({in0[59:56], in1[59:58]}, pp478);
level0_mult lvl0_mult479({in0[63:60], in1[59:58]}, pp479);
level0_mult lvl0_mult480({in0[3:0], in1[61:60]}, pp480);
level0_mult lvl0_mult481({in0[7:4], in1[61:60]}, pp481);
level0_mult lvl0_mult482({in0[11:8], in1[61:60]}, pp482);
level0_mult lvl0_mult483({in0[15:12], in1[61:60]}, pp483);
level0_mult lvl0_mult484({in0[19:16], in1[61:60]}, pp484);
level0_mult lvl0_mult485({in0[23:20], in1[61:60]}, pp485);
level0_mult lvl0_mult486({in0[27:24], in1[61:60]}, pp486);
level0_mult lvl0_mult487({in0[31:28], in1[61:60]}, pp487);
level0_mult lvl0_mult488({in0[35:32], in1[61:60]}, pp488);
level0_mult lvl0_mult489({in0[39:36], in1[61:60]}, pp489);
level0_mult lvl0_mult490({in0[43:40], in1[61:60]}, pp490);
level0_mult lvl0_mult491({in0[47:44], in1[61:60]}, pp491);
level0_mult lvl0_mult492({in0[51:48], in1[61:60]}, pp492);
level0_mult lvl0_mult493({in0[55:52], in1[61:60]}, pp493);
level0_mult lvl0_mult494({in0[59:56], in1[61:60]}, pp494);
level0_mult lvl0_mult495({in0[63:60], in1[61:60]}, pp495);
level0_mult lvl0_mult496({in0[3:0], in1[63:62]}, pp496);
level0_mult lvl0_mult497({in0[7:4], in1[63:62]}, pp497);
level0_mult lvl0_mult498({in0[11:8], in1[63:62]}, pp498);
level0_mult lvl0_mult499({in0[15:12], in1[63:62]}, pp499);
level0_mult lvl0_mult500({in0[19:16], in1[63:62]}, pp500);
level0_mult lvl0_mult501({in0[23:20], in1[63:62]}, pp501);
level0_mult lvl0_mult502({in0[27:24], in1[63:62]}, pp502);
level0_mult lvl0_mult503({in0[31:28], in1[63:62]}, pp503);
level0_mult lvl0_mult504({in0[35:32], in1[63:62]}, pp504);
level0_mult lvl0_mult505({in0[39:36], in1[63:62]}, pp505);
level0_mult lvl0_mult506({in0[43:40], in1[63:62]}, pp506);
level0_mult lvl0_mult507({in0[47:44], in1[63:62]}, pp507);
level0_mult lvl0_mult508({in0[51:48], in1[63:62]}, pp508);
level0_mult lvl0_mult509({in0[55:52], in1[63:62]}, pp509);
level0_mult lvl0_mult510({in0[59:56], in1[63:62]}, pp510);
level0_mult lvl0_mult511({in0[63:60], in1[63:62]}, pp511);


// level 0
wire [2:0]  gpcOutL0_0;
wire [2:0]  gpcOutL0_1;
wire [2:0]  gpcOutL0_2;
wire [2:0]  gpcOutL0_3;
wire [2:0]  gpcOutL0_4;
wire [2:0]  gpcOutL0_5;
wire [2:0]  gpcOutL0_6;
wire [2:0]  gpcOutL0_7;
wire [2:0]  gpcOutL0_8;
wire [2:0]  gpcOutL0_9;
wire [2:0]  gpcOutL0_10;
wire [2:0]  gpcOutL0_11;
wire [2:0]  gpcOutL0_12;
wire [2:0]  gpcOutL0_13;
wire [2:0]  gpcOutL0_14;
wire [2:0]  gpcOutL0_15;
wire [2:0]  gpcOutL0_16;
wire [2:0]  gpcOutL0_17;
wire [2:0]  gpcOutL0_18;
wire [2:0]  gpcOutL0_19;
wire [2:0]  gpcOutL0_20;
wire [2:0]  gpcOutL0_21;
wire [2:0]  gpcOutL0_22;
wire [2:0]  gpcOutL0_23;
wire [2:0]  gpcOutL0_24;
wire [2:0]  gpcOutL0_25;
wire [2:0]  gpcOutL0_26;
wire [2:0]  gpcOutL0_27;
wire [2:0]  gpcOutL0_28;
wire [2:0]  gpcOutL0_29;
wire [2:0]  gpcOutL0_30;
wire [2:0]  gpcOutL0_31;
wire [2:0]  gpcOutL0_32;
wire [2:0]  gpcOutL0_33;
wire [2:0]  gpcOutL0_34;
wire [2:0]  gpcOutL0_35;
wire [2:0]  gpcOutL0_36;
wire [2:0]  gpcOutL0_37;
wire [2:0]  gpcOutL0_38;
wire [2:0]  gpcOutL0_39;
wire [2:0]  gpcOutL0_40;
wire [2:0]  gpcOutL0_41;
wire [2:0]  gpcOutL0_42;
wire [2:0]  gpcOutL0_43;
wire [2:0]  gpcOutL0_44;
wire [2:0]  gpcOutL0_45;
wire [2:0]  gpcOutL0_46;
wire [2:0]  gpcOutL0_47;
wire [2:0]  gpcOutL0_48;
wire [2:0]  gpcOutL0_49;
wire [2:0]  gpcOutL0_50;
wire [2:0]  gpcOutL0_51;
wire [2:0]  gpcOutL0_52;
wire [2:0]  gpcOutL0_53;
wire [2:0]  gpcOutL0_54;
wire [2:0]  gpcOutL0_55;
wire [2:0]  gpcOutL0_56;
wire [2:0]  gpcOutL0_57;
wire [2:0]  gpcOutL0_58;
wire [2:0]  gpcOutL0_59;
wire [2:0]  gpcOutL0_60;
wire [2:0]  gpcOutL0_61;
wire [2:0]  gpcOutL0_62;
wire [2:0]  gpcOutL0_63;
wire [2:0]  gpcOutL0_64;
wire [2:0]  gpcOutL0_65;
wire [2:0]  gpcOutL0_66;
wire [2:0]  gpcOutL0_67;
wire [2:0]  gpcOutL0_68;
wire [2:0]  gpcOutL0_69;
wire [2:0]  gpcOutL0_70;
wire [2:0]  gpcOutL0_71;
wire [2:0]  gpcOutL0_72;
wire [2:0]  gpcOutL0_73;
wire [2:0]  gpcOutL0_74;
wire [2:0]  gpcOutL0_75;
wire [2:0]  gpcOutL0_76;
wire [2:0]  gpcOutL0_77;
wire [2:0]  gpcOutL0_78;
wire [2:0]  gpcOutL0_79;
wire [2:0]  gpcOutL0_80;
wire [2:0]  gpcOutL0_81;
wire [2:0]  gpcOutL0_82;
wire [2:0]  gpcOutL0_83;
wire [2:0]  gpcOutL0_84;
wire [2:0]  gpcOutL0_85;
wire [2:0]  gpcOutL0_86;
wire [2:0]  gpcOutL0_87;
wire [2:0]  gpcOutL0_88;
wire [2:0]  gpcOutL0_89;
wire [2:0]  gpcOutL0_90;
wire [2:0]  gpcOutL0_91;
wire [2:0]  gpcOutL0_92;
wire [2:0]  gpcOutL0_93;
wire [2:0]  gpcOutL0_94;
wire [2:0]  gpcOutL0_95;
wire [2:0]  gpcOutL0_96;
wire [2:0]  gpcOutL0_97;
wire [2:0]  gpcOutL0_98;
wire [2:0]  gpcOutL0_99;
wire [2:0]  gpcOutL0_100;
wire [2:0]  gpcOutL0_101;
wire [2:0]  gpcOutL0_102;
wire [2:0]  gpcOutL0_103;
wire [2:0]  gpcOutL0_104;
wire [2:0]  gpcOutL0_105;
wire [2:0]  gpcOutL0_106;
wire [2:0]  gpcOutL0_107;
wire [2:0]  gpcOutL0_108;
wire [2:0]  gpcOutL0_109;
wire [2:0]  gpcOutL0_110;
wire [2:0]  gpcOutL0_111;
wire [2:0]  gpcOutL0_112;
wire [2:0]  gpcOutL0_113;
wire [2:0]  gpcOutL0_114;
wire [2:0]  gpcOutL0_115;
wire [2:0]  gpcOutL0_116;
wire [2:0]  gpcOutL0_117;
wire [2:0]  gpcOutL0_118;
wire [2:0]  gpcOutL0_119;
wire [2:0]  gpcOutL0_120;
wire [2:0]  gpcOutL0_121;
wire [2:0]  gpcOutL0_122;
wire [2:0]  gpcOutL0_123;
wire [2:0]  gpcOutL0_124;
wire [2:0]  gpcOutL0_125;
wire [2:0]  gpcOutL0_126;
wire [2:0]  gpcOutL0_127;
wire [2:0]  gpcOutL0_128;
wire [2:0]  gpcOutL0_129;
wire [2:0]  gpcOutL0_130;
wire [2:0]  gpcOutL0_131;
wire [2:0]  gpcOutL0_132;
wire [2:0]  gpcOutL0_133;
wire [2:0]  gpcOutL0_134;
wire [2:0]  gpcOutL0_135;
wire [2:0]  gpcOutL0_136;
wire [2:0]  gpcOutL0_137;
wire [2:0]  gpcOutL0_138;
wire [2:0]  gpcOutL0_139;
wire [2:0]  gpcOutL0_140;
wire [2:0]  gpcOutL0_141;
wire [2:0]  gpcOutL0_142;
wire [2:0]  gpcOutL0_143;
wire [2:0]  gpcOutL0_144;
wire [2:0]  gpcOutL0_145;
wire [2:0]  gpcOutL0_146;
wire [2:0]  gpcOutL0_147;
wire [2:0]  gpcOutL0_148;
wire [2:0]  gpcOutL0_149;
wire [2:0]  gpcOutL0_150;
wire [2:0]  gpcOutL0_151;
wire [2:0]  gpcOutL0_152;
wire [2:0]  gpcOutL0_153;
wire [2:0]  gpcOutL0_154;
wire [2:0]  gpcOutL0_155;
wire [2:0]  gpcOutL0_156;
wire [2:0]  gpcOutL0_157;
wire [2:0]  gpcOutL0_158;
wire [2:0]  gpcOutL0_159;
wire [2:0]  gpcOutL0_160;
wire [2:0]  gpcOutL0_161;
wire [2:0]  gpcOutL0_162;
wire [2:0]  gpcOutL0_163;
wire [2:0]  gpcOutL0_164;
wire [2:0]  gpcOutL0_165;
wire [2:0]  gpcOutL0_166;
wire [2:0]  gpcOutL0_167;
wire [2:0]  gpcOutL0_168;
wire [2:0]  gpcOutL0_169;
wire [2:0]  gpcOutL0_170;
wire [2:0]  gpcOutL0_171;
wire [2:0]  gpcOutL0_172;
wire [2:0]  gpcOutL0_173;
wire [2:0]  gpcOutL0_174;
wire [2:0]  gpcOutL0_175;
wire [2:0]  gpcOutL0_176;
wire [2:0]  gpcOutL0_177;
wire [2:0]  gpcOutL0_178;
wire [2:0]  gpcOutL0_179;
wire [2:0]  gpcOutL0_180;
wire [2:0]  gpcOutL0_181;
wire [2:0]  gpcOutL0_182;
wire [2:0]  gpcOutL0_183;
wire [2:0]  gpcOutL0_184;
wire [2:0]  gpcOutL0_185;
wire [2:0]  gpcOutL0_186;
wire [2:0]  gpcOutL0_187;
wire [2:0]  gpcOutL0_188;
wire [2:0]  gpcOutL0_189;
wire [2:0]  gpcOutL0_190;
wire [2:0]  gpcOutL0_191;
wire [2:0]  gpcOutL0_192;
wire [2:0]  gpcOutL0_193;
wire [2:0]  gpcOutL0_194;
wire [2:0]  gpcOutL0_195;
wire [2:0]  gpcOutL0_196;
wire [2:0]  gpcOutL0_197;
wire [2:0]  gpcOutL0_198;
wire [2:0]  gpcOutL0_199;
wire [2:0]  gpcOutL0_200;
wire [2:0]  gpcOutL0_201;
wire [2:0]  gpcOutL0_202;
wire [2:0]  gpcOutL0_203;
wire [2:0]  gpcOutL0_204;
wire [2:0]  gpcOutL0_205;
wire [2:0]  gpcOutL0_206;
wire [2:0]  gpcOutL0_207;
wire [2:0]  gpcOutL0_208;
wire [2:0]  gpcOutL0_209;
wire [2:0]  gpcOutL0_210;
wire [2:0]  gpcOutL0_211;
wire [2:0]  gpcOutL0_212;
wire [2:0]  gpcOutL0_213;
wire [2:0]  gpcOutL0_214;
wire [2:0]  gpcOutL0_215;
wire [2:0]  gpcOutL0_216;
wire [2:0]  gpcOutL0_217;
wire [2:0]  gpcOutL0_218;
wire [2:0]  gpcOutL0_219;
wire [2:0]  gpcOutL0_220;
wire [2:0]  gpcOutL0_221;
wire [2:0]  gpcOutL0_222;
wire [2:0]  gpcOutL0_223;
wire [2:0]  gpcOutL0_224;
wire [2:0]  gpcOutL0_225;
wire [2:0]  gpcOutL0_226;
wire [2:0]  gpcOutL0_227;
wire [2:0]  gpcOutL0_228;
wire [2:0]  gpcOutL0_229;
wire [2:0]  gpcOutL0_230;
wire [2:0]  gpcOutL0_231;
wire [2:0]  gpcOutL0_232;
wire [2:0]  gpcOutL0_233;
wire [2:0]  gpcOutL0_234;
wire [2:0]  gpcOutL0_235;
wire [2:0]  gpcOutL0_236;
wire [2:0]  gpcOutL0_237;
wire [2:0]  gpcOutL0_238;
wire [2:0]  gpcOutL0_239;
wire [2:0]  gpcOutL0_240;
wire [2:0]  gpcOutL0_241;
wire [2:0]  gpcOutL0_242;
wire [2:0]  gpcOutL0_243;
wire [2:0]  gpcOutL0_244;
wire [2:0]  gpcOutL0_245;
wire [2:0]  gpcOutL0_246;
wire [2:0]  gpcOutL0_247;
wire [2:0]  gpcOutL0_248;
wire [2:0]  gpcOutL0_249;
wire [2:0]  gpcOutL0_250;
wire [2:0]  gpcOutL0_251;
wire [2:0]  gpcOutL0_252;
wire [2:0]  gpcOutL0_253;
wire [2:0]  gpcOutL0_254;
wire [2:0]  gpcOutL0_255;
wire [2:0]  gpcOutL0_256;
wire [2:0]  gpcOutL0_257;
wire [2:0]  gpcOutL0_258;
wire [2:0]  gpcOutL0_259;
wire [2:0]  gpcOutL0_260;
wire [2:0]  gpcOutL0_261;
wire [2:0]  gpcOutL0_262;
wire [2:0]  gpcOutL0_263;
wire [2:0]  gpcOutL0_264;
wire [2:0]  gpcOutL0_265;
wire [2:0]  gpcOutL0_266;
wire [2:0]  gpcOutL0_267;
wire [2:0]  gpcOutL0_268;
wire [2:0]  gpcOutL0_269;
wire [2:0]  gpcOutL0_270;
wire [2:0]  gpcOutL0_271;
wire [2:0]  gpcOutL0_272;
wire [2:0]  gpcOutL0_273;
wire [2:0]  gpcOutL0_274;
wire [2:0]  gpcOutL0_275;
wire [2:0]  gpcOutL0_276;
wire [2:0]  gpcOutL0_277;
wire [2:0]  gpcOutL0_278;
wire [2:0]  gpcOutL0_279;
wire [2:0]  gpcOutL0_280;
wire [2:0]  gpcOutL0_281;
wire [2:0]  gpcOutL0_282;
wire [2:0]  gpcOutL0_283;
wire [2:0]  gpcOutL0_284;
wire [2:0]  gpcOutL0_285;
wire [2:0]  gpcOutL0_286;
wire [2:0]  gpcOutL0_287;
wire [2:0]  gpcOutL0_288;
wire [2:0]  gpcOutL0_289;
wire [2:0]  gpcOutL0_290;
wire [2:0]  gpcOutL0_291;
wire [2:0]  gpcOutL0_292;
wire [2:0]  gpcOutL0_293;
wire [2:0]  gpcOutL0_294;
wire [2:0]  gpcOutL0_295;
wire [2:0]  gpcOutL0_296;
wire [2:0]  gpcOutL0_297;
wire [2:0]  gpcOutL0_298;
wire [2:0]  gpcOutL0_299;
wire [2:0]  gpcOutL0_300;
wire [2:0]  gpcOutL0_301;
wire [2:0]  gpcOutL0_302;
wire [2:0]  gpcOutL0_303;
wire [2:0]  gpcOutL0_304;
wire [2:0]  gpcOutL0_305;
wire [2:0]  gpcOutL0_306;
wire [2:0]  gpcOutL0_307;
wire [2:0]  gpcOutL0_308;
wire [2:0]  gpcOutL0_309;
wire [2:0]  gpcOutL0_310;
wire [2:0]  gpcOutL0_311;
wire [2:0]  gpcOutL0_312;
wire [2:0]  gpcOutL0_313;
wire [2:0]  gpcOutL0_314;
wire [2:0]  gpcOutL0_315;
wire [2:0]  gpcOutL0_316;
wire [2:0]  gpcOutL0_317;
wire [2:0]  gpcOutL0_318;
wire [2:0]  gpcOutL0_319;
wire [2:0]  gpcOutL0_320;
wire [2:0]  gpcOutL0_321;
wire [2:0]  gpcOutL0_322;
wire [2:0]  gpcOutL0_323;
wire [2:0]  gpcOutL0_324;
wire [2:0]  gpcOutL0_325;
wire [2:0]  gpcOutL0_326;
wire [2:0]  gpcOutL0_327;
wire [2:0]  gpcOutL0_328;
wire [2:0]  gpcOutL0_329;
wire [2:0]  gpcOutL0_330;
wire [2:0]  gpcOutL0_331;
wire [2:0]  gpcOutL0_332;
wire [2:0]  gpcOutL0_333;
wire [2:0]  gpcOutL0_334;
wire [2:0]  gpcOutL0_335;
wire [2:0]  gpcOutL0_336;
wire [2:0]  gpcOutL0_337;
wire [2:0]  gpcOutL0_338;
wire [2:0]  gpcOutL0_339;
wire [2:0]  gpcOutL0_340;
wire [2:0]  gpcOutL0_341;
wire [2:0]  gpcOutL0_342;
wire [2:0]  gpcOutL0_343;
wire [2:0]  gpcOutL0_344;
wire [2:0]  gpcOutL0_345;
wire [2:0]  gpcOutL0_346;
wire [2:0]  gpcOutL0_347;
wire [2:0]  gpcOutL0_348;
wire [2:0]  gpcOutL0_349;
wire [2:0]  gpcOutL0_350;
wire [2:0]  gpcOutL0_351;
wire [2:0]  gpcOutL0_352;
wire [2:0]  gpcOutL0_353;
wire [2:0]  gpcOutL0_354;
wire [2:0]  gpcOutL0_355;
wire [2:0]  gpcOutL0_356;
wire [2:0]  gpcOutL0_357;
wire [2:0]  gpcOutL0_358;
wire [2:0]  gpcOutL0_359;
wire [2:0]  gpcOutL0_360;
wire [2:0]  gpcOutL0_361;
wire [2:0]  gpcOutL0_362;
wire [2:0]  gpcOutL0_363;
wire [2:0]  gpcOutL0_364;
wire [2:0]  gpcOutL0_365;
wire [2:0]  gpcOutL0_366;
wire [2:0]  gpcOutL0_367;
wire [2:0]  gpcOutL0_368;
wire [2:0]  gpcOutL0_369;
wire [2:0]  gpcOutL0_370;
wire [2:0]  gpcOutL0_371;
wire [2:0]  gpcOutL0_372;
wire [2:0]  gpcOutL0_373;
wire [2:0]  gpcOutL0_374;
wire [2:0]  gpcOutL0_375;
wire [2:0]  gpcOutL0_376;
wire [2:0]  gpcOutL0_377;
wire [2:0]  gpcOutL0_378;
wire [2:0]  gpcOutL0_379;
wire [2:0]  gpcOutL0_380;
wire [2:0]  gpcOutL0_381;
wire [2:0]  gpcOutL0_382;
wire [2:0]  gpcOutL0_383;
wire [2:0]  gpcOutL0_384;
wire [2:0]  gpcOutL0_385;
wire [2:0]  gpcOutL0_386;
wire [2:0]  gpcOutL0_387;
wire [2:0]  gpcOutL0_388;
wire [2:0]  gpcOutL0_389;
wire [2:0]  gpcOutL0_390;
wire [2:0]  gpcOutL0_391;
wire [2:0]  gpcOutL0_392;
wire [2:0]  gpcOutL0_393;
wire [2:0]  gpcOutL0_394;
wire [2:0]  gpcOutL0_395;
wire [2:0]  gpcOutL0_396;
wire [2:0]  gpcOutL0_397;
wire [2:0]  gpcOutL0_398;
wire [2:0]  gpcOutL0_399;
wire [2:0]  gpcOutL0_400;
wire [2:0]  gpcOutL0_401;
wire [2:0]  gpcOutL0_402;
wire [2:0]  gpcOutL0_403;
wire [2:0]  gpcOutL0_404;
wire [2:0]  gpcOutL0_405;
wire [2:0]  gpcOutL0_406;
wire [2:0]  gpcOutL0_407;
wire [2:0]  gpcOutL0_408;
wire [2:0]  gpcOutL0_409;
wire [2:0]  gpcOutL0_410;
wire [2:0]  gpcOutL0_411;
wire [2:0]  gpcOutL0_412;
wire [2:0]  gpcOutL0_413;
wire [2:0]  gpcOutL0_414;
wire [2:0]  gpcOutL0_415;
wire [2:0]  gpcOutL0_416;
wire [2:0]  gpcOutL0_417;
wire [2:0]  gpcOutL0_418;
wire [2:0]  gpcOutL0_419;
wire [2:0]  gpcOutL0_420;
wire [2:0]  gpcOutL0_421;
wire [2:0]  gpcOutL0_422;
wire [2:0]  gpcOutL0_423;
wire [2:0]  gpcOutL0_424;
wire [2:0]  gpcOutL0_425;
wire [2:0]  gpcOutL0_426;
wire [2:0]  gpcOutL0_427;
wire [2:0]  gpcOutL0_428;
wire [2:0]  gpcOutL0_429;
wire [2:0]  gpcOutL0_430;
wire [2:0]  gpcOutL0_431;
wire [2:0]  gpcOutL0_432;
wire [2:0]  gpcOutL0_433;
wire [2:0]  gpcOutL0_434;
wire [2:0]  gpcOutL0_435;
wire [2:0]  gpcOutL0_436;
wire [2:0]  gpcOutL0_437;
wire [2:0]  gpcOutL0_438;
wire [2:0]  gpcOutL0_439;
wire [2:0]  gpcOutL0_440;
wire [2:0]  gpcOutL0_441;
wire [2:0]  gpcOutL0_442;
wire [2:0]  gpcOutL0_443;
wire [2:0]  gpcOutL0_444;
wire [2:0]  gpcOutL0_445;
wire [2:0]  gpcOutL0_446;
wire [2:0]  gpcOutL0_447;
wire [2:0]  gpcOutL0_448;
wire [2:0]  gpcOutL0_449;
wire [2:0]  gpcOutL0_450;
wire [2:0]  gpcOutL0_451;
wire [2:0]  gpcOutL0_452;
wire [2:0]  gpcOutL0_453;
wire [2:0]  gpcOutL0_454;
wire [2:0]  gpcOutL0_455;
wire [2:0]  gpcOutL0_456;
wire [2:0]  gpcOutL0_457;
wire [2:0]  gpcOutL0_458;
wire [2:0]  gpcOutL0_459;
wire [2:0]  gpcOutL0_460;
wire [2:0]  gpcOutL0_461;
wire [2:0]  gpcOutL0_462;
wire [2:0]  gpcOutL0_463;
wire [2:0]  gpcOutL0_464;
wire [2:0]  gpcOutL0_465;
wire [2:0]  gpcOutL0_466;
wire [2:0]  gpcOutL0_467;
wire [2:0]  gpcOutL0_468;
wire [2:0]  gpcOutL0_469;
wire [2:0]  gpcOutL0_470;
wire [2:0]  gpcOutL0_471;
wire [2:0]  gpcOutL0_472;
wire [2:0]  gpcOutL0_473;
wire [2:0]  gpcOutL0_474;
wire [2:0]  gpcOutL0_475;
wire [2:0]  gpcOutL0_476;
wire [2:0]  gpcOutL0_477;
wire [2:0]  gpcOutL0_478;
wire [2:0]  gpcOutL0_479;
wire [2:0]  gpcOutL0_480;
wire [2:0]  gpcOutL0_481;
wire [2:0]  gpcOutL0_482;
wire [2:0]  gpcOutL0_483;
wire [2:0]  gpcOutL0_484;
wire [2:0]  gpcOutL0_485;
wire [2:0]  gpcOutL0_486;
wire [2:0]  gpcOutL0_487;
wire [2:0]  gpcOutL0_488;
wire [2:0]  gpcOutL0_489;
wire [2:0]  gpcOutL0_490;
wire [2:0]  gpcOutL0_491;
wire [2:0]  gpcOutL0_492;
wire [2:0]  gpcOutL0_493;
wire [2:0]  gpcOutL0_494;
wire [1:0]  gpcOutL0_495;
wire [1:0]  gpcOutL0_496;
wire [1:0]  gpcOutL0_497;
wire [1:0]  gpcOutL0_498;
wire [1:0]  gpcOutL0_499;
wire [1:0]  gpcOutL0_500;
wire [1:0]  gpcOutL0_501;
wire [1:0]  gpcOutL0_502;
wire [1:0]  gpcOutL0_503;
wire [1:0]  gpcOutL0_504;
wire [1:0]  gpcOutL0_505;
wire [1:0]  gpcOutL0_506;
wire [1:0]  gpcOutL0_507;
wire [1:0]  gpcOutL0_508;
wire [1:0]  gpcOutL0_509;
wire [1:0]  gpcOutL0_510;
wire [1:0]  gpcOutL0_511;
wire [2:0]  gpcOutL0_512;
wire [2:0]  gpcOutL0_513;
wire [2:0]  gpcOutL0_514;
wire [2:0]  gpcOutL0_515;
wire [2:0]  gpcOutL0_516;
wire [2:0]  gpcOutL0_517;
wire [2:0]  gpcOutL0_518;
wire [2:0]  gpcOutL0_519;

gpc006 gpcL0_0 ({pp64[0], pp48[2], pp33[0], pp32[4], pp17[2], pp2[0]}, gpcOutL0_0);
gpc006 gpcL0_1 ({pp64[1], pp48[3], pp33[1], pp32[5], pp17[3], pp2[1]}, gpcOutL0_1);
gpc006 gpcL0_2 ({pp80[0], pp64[2], pp49[0], pp48[4], pp33[2], pp18[0]}, gpcOutL0_2);
gpc006 gpcL0_3 ({pp80[1], pp64[3], pp49[1], pp48[5], pp33[3], pp18[1]}, gpcOutL0_3);
gpc006 gpcL0_4 ({pp96[0], pp80[2], pp65[0], pp64[4], pp49[2], pp34[0]}, gpcOutL0_4);
gpc006 gpcL0_5 ({pp96[1], pp80[3], pp65[1], pp64[5], pp49[3], pp34[1]}, gpcOutL0_5);
gpc006 gpcL0_6 ({pp112[0], pp96[2], pp81[0], pp80[4], pp65[2], pp50[0]}, gpcOutL0_6);
gpc006 gpcL0_7 ({pp112[1], pp96[3], pp81[1], pp80[5], pp65[3], pp50[1]}, gpcOutL0_7);
gpc006 gpcL0_8 ({pp128[0], pp112[2], pp97[0], pp96[4], pp81[2], pp66[0]}, gpcOutL0_8);
gpc006 gpcL0_9 ({pp128[1], pp112[3], pp97[1], pp96[5], pp81[3], pp66[1]}, gpcOutL0_9);
gpc006 gpcL0_10 ({pp144[0], pp128[2], pp113[0], pp112[4], pp97[2], pp82[0]}, gpcOutL0_10);
gpc006 gpcL0_11 ({pp144[1], pp128[3], pp113[1], pp112[5], pp97[3], pp82[1]}, gpcOutL0_11);
gpc006 gpcL0_12 ({pp160[0], pp144[2], pp129[0], pp128[4], pp113[2], pp98[0]}, gpcOutL0_12);
gpc006 gpcL0_13 ({pp160[1], pp144[3], pp129[1], pp128[5], pp113[3], pp98[1]}, gpcOutL0_13);
gpc006 gpcL0_14 ({pp176[0], pp160[2], pp145[0], pp144[4], pp129[2], pp114[0]}, gpcOutL0_14);
gpc006 gpcL0_15 ({pp176[1], pp160[3], pp145[1], pp144[5], pp129[3], pp114[1]}, gpcOutL0_15);
gpc006 gpcL0_16 ({pp192[0], pp176[2], pp161[0], pp160[4], pp145[2], pp130[0]}, gpcOutL0_16);
gpc006 gpcL0_17 ({pp192[1], pp176[3], pp161[1], pp160[5], pp145[3], pp130[1]}, gpcOutL0_17);
gpc006 gpcL0_18 ({pp208[0], pp192[2], pp177[0], pp176[4], pp161[2], pp146[0]}, gpcOutL0_18);
gpc006 gpcL0_19 ({pp208[1], pp192[3], pp177[1], pp176[5], pp161[3], pp146[1]}, gpcOutL0_19);
gpc006 gpcL0_20 ({pp224[0], pp208[2], pp193[0], pp192[4], pp177[2], pp162[0]}, gpcOutL0_20);
gpc006 gpcL0_21 ({pp224[1], pp208[3], pp193[1], pp192[5], pp177[3], pp162[1]}, gpcOutL0_21);
gpc006 gpcL0_22 ({pp240[0], pp224[2], pp209[0], pp208[4], pp193[2], pp178[0]}, gpcOutL0_22);
gpc006 gpcL0_23 ({pp240[1], pp224[3], pp209[1], pp208[5], pp193[3], pp178[1]}, gpcOutL0_23);
gpc006 gpcL0_24 ({pp256[0], pp240[2], pp225[0], pp224[4], pp209[2], pp194[0]}, gpcOutL0_24);
gpc006 gpcL0_25 ({pp256[1], pp240[3], pp225[1], pp224[5], pp209[3], pp194[1]}, gpcOutL0_25);
gpc006 gpcL0_26 ({pp272[0], pp256[2], pp241[0], pp240[4], pp225[2], pp210[0]}, gpcOutL0_26);
gpc006 gpcL0_27 ({pp272[1], pp256[3], pp241[1], pp240[5], pp225[3], pp210[1]}, gpcOutL0_27);
gpc006 gpcL0_28 ({pp288[0], pp272[2], pp257[0], pp256[4], pp241[2], pp226[0]}, gpcOutL0_28);
gpc006 gpcL0_29 ({pp288[1], pp272[3], pp257[1], pp256[5], pp241[3], pp226[1]}, gpcOutL0_29);
gpc006 gpcL0_30 ({pp304[0], pp288[2], pp273[0], pp272[4], pp257[2], pp242[0]}, gpcOutL0_30);
gpc006 gpcL0_31 ({pp304[1], pp288[3], pp273[1], pp272[5], pp257[3], pp242[1]}, gpcOutL0_31);
gpc006 gpcL0_32 ({pp320[0], pp304[2], pp289[0], pp288[4], pp273[2], pp258[0]}, gpcOutL0_32);
gpc006 gpcL0_33 ({pp320[1], pp304[3], pp289[1], pp288[5], pp273[3], pp258[1]}, gpcOutL0_33);
gpc006 gpcL0_34 ({pp336[0], pp320[2], pp305[0], pp304[4], pp289[2], pp274[0]}, gpcOutL0_34);
gpc006 gpcL0_35 ({pp336[1], pp320[3], pp305[1], pp304[5], pp289[3], pp274[1]}, gpcOutL0_35);
gpc006 gpcL0_36 ({pp352[0], pp336[2], pp321[0], pp320[4], pp305[2], pp290[0]}, gpcOutL0_36);
gpc006 gpcL0_37 ({pp352[1], pp336[3], pp321[1], pp320[5], pp305[3], pp290[1]}, gpcOutL0_37);
gpc006 gpcL0_38 ({pp368[0], pp352[2], pp337[0], pp336[4], pp321[2], pp306[0]}, gpcOutL0_38);
gpc006 gpcL0_39 ({pp368[1], pp352[3], pp337[1], pp336[5], pp321[3], pp306[1]}, gpcOutL0_39);
gpc006 gpcL0_40 ({pp384[0], pp368[2], pp353[0], pp352[4], pp337[2], pp322[0]}, gpcOutL0_40);
gpc006 gpcL0_41 ({pp384[1], pp368[3], pp353[1], pp352[5], pp337[3], pp322[1]}, gpcOutL0_41);
gpc006 gpcL0_42 ({pp400[0], pp384[2], pp369[0], pp368[4], pp353[2], pp338[0]}, gpcOutL0_42);
gpc006 gpcL0_43 ({pp400[1], pp384[3], pp369[1], pp368[5], pp353[3], pp338[1]}, gpcOutL0_43);
gpc006 gpcL0_44 ({pp416[0], pp400[2], pp385[0], pp384[4], pp369[2], pp354[0]}, gpcOutL0_44);
gpc006 gpcL0_45 ({pp416[1], pp400[3], pp385[1], pp384[5], pp369[3], pp354[1]}, gpcOutL0_45);
gpc006 gpcL0_46 ({pp432[0], pp416[2], pp401[0], pp400[4], pp385[2], pp370[0]}, gpcOutL0_46);
gpc006 gpcL0_47 ({pp432[1], pp416[3], pp401[1], pp400[5], pp385[3], pp370[1]}, gpcOutL0_47);
gpc006 gpcL0_48 ({pp448[0], pp432[2], pp417[0], pp416[4], pp401[2], pp386[0]}, gpcOutL0_48);
gpc006 gpcL0_49 ({pp448[1], pp432[3], pp417[1], pp416[5], pp401[3], pp386[1]}, gpcOutL0_49);
gpc006 gpcL0_50 ({pp464[0], pp448[2], pp433[0], pp432[4], pp417[2], pp402[0]}, gpcOutL0_50);
gpc006 gpcL0_51 ({pp464[1], pp448[3], pp433[1], pp432[5], pp417[3], pp402[1]}, gpcOutL0_51);
gpc006 gpcL0_52 ({pp480[0], pp464[2], pp449[0], pp448[4], pp433[2], pp418[0]}, gpcOutL0_52);
gpc006 gpcL0_53 ({pp480[1], pp464[3], pp449[1], pp448[5], pp433[3], pp418[1]}, gpcOutL0_53);
gpc006 gpcL0_54 ({pp496[0], pp480[2], pp465[0], pp464[4], pp449[2], pp434[0]}, gpcOutL0_54);
gpc006 gpcL0_55 ({pp496[1], pp480[3], pp465[1], pp464[5], pp449[3], pp434[1]}, gpcOutL0_55);
gpc006 gpcL0_56 ({pp496[2], pp481[0], pp480[4], pp465[2], pp450[0], pp449[4]}, gpcOutL0_56);
gpc006 gpcL0_57 ({pp496[3], pp481[1], pp480[5], pp465[3], pp450[1], pp449[5]}, gpcOutL0_57);
gpc006 gpcL0_58 ({pp497[0], pp496[4], pp481[2], pp466[0], pp465[4], pp450[2]}, gpcOutL0_58);
gpc006 gpcL0_59 ({pp497[1], pp496[5], pp481[3], pp466[1], pp465[5], pp450[3]}, gpcOutL0_59);
gpc006 gpcL0_60 ({pp497[2], pp482[0], pp481[4], pp466[2], pp451[0], pp450[4]}, gpcOutL0_60);
gpc006 gpcL0_61 ({pp497[3], pp482[1], pp481[5], pp466[3], pp451[1], pp450[5]}, gpcOutL0_61);
gpc006 gpcL0_62 ({pp498[0], pp497[4], pp482[2], pp467[0], pp466[4], pp451[2]}, gpcOutL0_62);
gpc006 gpcL0_63 ({pp498[1], pp497[5], pp482[3], pp467[1], pp466[5], pp451[3]}, gpcOutL0_63);
gpc006 gpcL0_64 ({pp498[2], pp483[0], pp482[4], pp467[2], pp452[0], pp451[4]}, gpcOutL0_64);
gpc006 gpcL0_65 ({pp498[3], pp483[1], pp482[5], pp467[3], pp452[1], pp451[5]}, gpcOutL0_65);
gpc006 gpcL0_66 ({pp499[0], pp498[4], pp483[2], pp468[0], pp467[4], pp452[2]}, gpcOutL0_66);
gpc006 gpcL0_67 ({pp499[1], pp498[5], pp483[3], pp468[1], pp467[5], pp452[3]}, gpcOutL0_67);
gpc006 gpcL0_68 ({pp499[2], pp484[0], pp483[4], pp468[2], pp453[0], pp452[4]}, gpcOutL0_68);
gpc006 gpcL0_69 ({pp499[3], pp484[1], pp483[5], pp468[3], pp453[1], pp452[5]}, gpcOutL0_69);
gpc006 gpcL0_70 ({pp500[0], pp499[4], pp484[2], pp469[0], pp468[4], pp453[2]}, gpcOutL0_70);
gpc006 gpcL0_71 ({pp500[1], pp499[5], pp484[3], pp469[1], pp468[5], pp453[3]}, gpcOutL0_71);
gpc006 gpcL0_72 ({pp500[2], pp485[0], pp484[4], pp469[2], pp454[0], pp453[4]}, gpcOutL0_72);
gpc006 gpcL0_73 ({pp500[3], pp485[1], pp484[5], pp469[3], pp454[1], pp453[5]}, gpcOutL0_73);
gpc006 gpcL0_74 ({pp501[0], pp500[4], pp485[2], pp470[0], pp469[4], pp454[2]}, gpcOutL0_74);
gpc006 gpcL0_75 ({pp501[1], pp500[5], pp485[3], pp470[1], pp469[5], pp454[3]}, gpcOutL0_75);
gpc006 gpcL0_76 ({pp501[2], pp486[0], pp485[4], pp470[2], pp455[0], pp454[4]}, gpcOutL0_76);
gpc006 gpcL0_77 ({pp501[3], pp486[1], pp485[5], pp470[3], pp455[1], pp454[5]}, gpcOutL0_77);
gpc006 gpcL0_78 ({pp502[0], pp501[4], pp486[2], pp471[0], pp470[4], pp455[2]}, gpcOutL0_78);
gpc006 gpcL0_79 ({pp502[1], pp501[5], pp486[3], pp471[1], pp470[5], pp455[3]}, gpcOutL0_79);
gpc006 gpcL0_80 ({pp502[2], pp487[0], pp486[4], pp471[2], pp456[0], pp455[4]}, gpcOutL0_80);
gpc006 gpcL0_81 ({pp502[3], pp487[1], pp486[5], pp471[3], pp456[1], pp455[5]}, gpcOutL0_81);
gpc006 gpcL0_82 ({pp503[0], pp502[4], pp487[2], pp472[0], pp471[4], pp456[2]}, gpcOutL0_82);
gpc006 gpcL0_83 ({pp503[1], pp502[5], pp487[3], pp472[1], pp471[5], pp456[3]}, gpcOutL0_83);
gpc006 gpcL0_84 ({pp503[2], pp488[0], pp487[4], pp472[2], pp457[0], pp456[4]}, gpcOutL0_84);
gpc006 gpcL0_85 ({pp503[3], pp488[1], pp487[5], pp472[3], pp457[1], pp456[5]}, gpcOutL0_85);
gpc006 gpcL0_86 ({pp504[0], pp503[4], pp488[2], pp473[0], pp472[4], pp457[2]}, gpcOutL0_86);
gpc006 gpcL0_87 ({pp504[1], pp503[5], pp488[3], pp473[1], pp472[5], pp457[3]}, gpcOutL0_87);
gpc006 gpcL0_88 ({pp504[2], pp489[0], pp488[4], pp473[2], pp458[0], pp457[4]}, gpcOutL0_88);
gpc006 gpcL0_89 ({pp504[3], pp489[1], pp488[5], pp473[3], pp458[1], pp457[5]}, gpcOutL0_89);
gpc006 gpcL0_90 ({pp505[0], pp504[4], pp489[2], pp474[0], pp473[4], pp458[2]}, gpcOutL0_90);
gpc006 gpcL0_91 ({pp505[1], pp504[5], pp489[3], pp474[1], pp473[5], pp458[3]}, gpcOutL0_91);
gpc006 gpcL0_92 ({pp505[2], pp490[0], pp489[4], pp474[2], pp459[0], pp458[4]}, gpcOutL0_92);
gpc006 gpcL0_93 ({pp505[3], pp490[1], pp489[5], pp474[3], pp459[1], pp458[5]}, gpcOutL0_93);
gpc006 gpcL0_94 ({pp506[0], pp505[4], pp490[2], pp475[0], pp474[4], pp459[2]}, gpcOutL0_94);
gpc006 gpcL0_95 ({pp506[1], pp505[5], pp490[3], pp475[1], pp474[5], pp459[3]}, gpcOutL0_95);
gpc006 gpcL0_96 ({pp506[2], pp491[0], pp490[4], pp475[2], pp460[0], pp459[4]}, gpcOutL0_96);
gpc006 gpcL0_97 ({pp506[3], pp491[1], pp490[5], pp475[3], pp460[1], pp459[5]}, gpcOutL0_97);
gpc006 gpcL0_98 ({pp507[0], pp506[4], pp491[2], pp476[0], pp475[4], pp460[2]}, gpcOutL0_98);
gpc006 gpcL0_99 ({pp507[1], pp506[5], pp491[3], pp476[1], pp475[5], pp460[3]}, gpcOutL0_99);
gpc006 gpcL0_100 ({pp507[2], pp492[0], pp491[4], pp476[2], pp461[0], pp460[4]}, gpcOutL0_100);
gpc006 gpcL0_101 ({pp507[3], pp492[1], pp491[5], pp476[3], pp461[1], pp460[5]}, gpcOutL0_101);
gpc006 gpcL0_102 ({pp508[0], pp507[4], pp492[2], pp477[0], pp476[4], pp461[2]}, gpcOutL0_102);
gpc006 gpcL0_103 ({pp508[1], pp507[5], pp492[3], pp477[1], pp476[5], pp461[3]}, gpcOutL0_103);
gpc006 gpcL0_104 ({pp508[2], pp493[0], pp492[4], pp477[2], pp462[0], pp461[4]}, gpcOutL0_104);
gpc006 gpcL0_105 ({pp508[3], pp493[1], pp492[5], pp477[3], pp462[1], pp461[5]}, gpcOutL0_105);
gpc006 gpcL0_106 ({pp509[0], pp508[4], pp493[2], pp478[0], pp477[4], pp462[2]}, gpcOutL0_106);
gpc006 gpcL0_107 ({pp509[1], pp508[5], pp493[3], pp478[1], pp477[5], pp462[3]}, gpcOutL0_107);
gpc006 gpcL0_108 ({pp509[2], pp494[0], pp493[4], pp478[2], pp463[0], pp462[4]}, gpcOutL0_108);
gpc006 gpcL0_109 ({pp509[3], pp494[1], pp493[5], pp478[3], pp463[1], pp462[5]}, gpcOutL0_109);
gpc006 gpcL0_110 ({pp510[0], pp509[4], pp494[2], pp479[0], pp478[4], pp463[2]}, gpcOutL0_110);
gpc006 gpcL0_111 ({pp510[1], pp509[5], pp494[3], pp479[1], pp478[5], pp463[3]}, gpcOutL0_111);
gpc006 gpcL0_112 ({pp65[4], pp50[2], pp35[0], pp34[4], pp19[2], pp4[0]}, gpcOutL0_112);
gpc006 gpcL0_113 ({pp65[5], pp50[3], pp35[1], pp34[5], pp19[3], pp4[1]}, gpcOutL0_113);
gpc006 gpcL0_114 ({pp81[4], pp66[2], pp51[0], pp50[4], pp35[2], pp20[0]}, gpcOutL0_114);
gpc006 gpcL0_115 ({pp81[5], pp66[3], pp51[1], pp50[5], pp35[3], pp20[1]}, gpcOutL0_115);
gpc006 gpcL0_116 ({pp97[4], pp82[2], pp67[0], pp66[4], pp51[2], pp36[0]}, gpcOutL0_116);
gpc006 gpcL0_117 ({pp97[5], pp82[3], pp67[1], pp66[5], pp51[3], pp36[1]}, gpcOutL0_117);
gpc006 gpcL0_118 ({pp113[4], pp98[2], pp83[0], pp82[4], pp67[2], pp52[0]}, gpcOutL0_118);
gpc006 gpcL0_119 ({pp113[5], pp98[3], pp83[1], pp82[5], pp67[3], pp52[1]}, gpcOutL0_119);
gpc006 gpcL0_120 ({pp129[4], pp114[2], pp99[0], pp98[4], pp83[2], pp68[0]}, gpcOutL0_120);
gpc006 gpcL0_121 ({pp129[5], pp114[3], pp99[1], pp98[5], pp83[3], pp68[1]}, gpcOutL0_121);
gpc006 gpcL0_122 ({pp145[4], pp130[2], pp115[0], pp114[4], pp99[2], pp84[0]}, gpcOutL0_122);
gpc006 gpcL0_123 ({pp145[5], pp130[3], pp115[1], pp114[5], pp99[3], pp84[1]}, gpcOutL0_123);
gpc006 gpcL0_124 ({pp161[4], pp146[2], pp131[0], pp130[4], pp115[2], pp100[0]}, gpcOutL0_124);
gpc006 gpcL0_125 ({pp161[5], pp146[3], pp131[1], pp130[5], pp115[3], pp100[1]}, gpcOutL0_125);
gpc006 gpcL0_126 ({pp177[4], pp162[2], pp147[0], pp146[4], pp131[2], pp116[0]}, gpcOutL0_126);
gpc006 gpcL0_127 ({pp177[5], pp162[3], pp147[1], pp146[5], pp131[3], pp116[1]}, gpcOutL0_127);
gpc006 gpcL0_128 ({pp193[4], pp178[2], pp163[0], pp162[4], pp147[2], pp132[0]}, gpcOutL0_128);
gpc006 gpcL0_129 ({pp193[5], pp178[3], pp163[1], pp162[5], pp147[3], pp132[1]}, gpcOutL0_129);
gpc006 gpcL0_130 ({pp209[4], pp194[2], pp179[0], pp178[4], pp163[2], pp148[0]}, gpcOutL0_130);
gpc006 gpcL0_131 ({pp209[5], pp194[3], pp179[1], pp178[5], pp163[3], pp148[1]}, gpcOutL0_131);
gpc006 gpcL0_132 ({pp225[4], pp210[2], pp195[0], pp194[4], pp179[2], pp164[0]}, gpcOutL0_132);
gpc006 gpcL0_133 ({pp225[5], pp210[3], pp195[1], pp194[5], pp179[3], pp164[1]}, gpcOutL0_133);
gpc006 gpcL0_134 ({pp241[4], pp226[2], pp211[0], pp210[4], pp195[2], pp180[0]}, gpcOutL0_134);
gpc006 gpcL0_135 ({pp241[5], pp226[3], pp211[1], pp210[5], pp195[3], pp180[1]}, gpcOutL0_135);
gpc006 gpcL0_136 ({pp257[4], pp242[2], pp227[0], pp226[4], pp211[2], pp196[0]}, gpcOutL0_136);
gpc006 gpcL0_137 ({pp257[5], pp242[3], pp227[1], pp226[5], pp211[3], pp196[1]}, gpcOutL0_137);
gpc006 gpcL0_138 ({pp273[4], pp258[2], pp243[0], pp242[4], pp227[2], pp212[0]}, gpcOutL0_138);
gpc006 gpcL0_139 ({pp273[5], pp258[3], pp243[1], pp242[5], pp227[3], pp212[1]}, gpcOutL0_139);
gpc006 gpcL0_140 ({pp289[4], pp274[2], pp259[0], pp258[4], pp243[2], pp228[0]}, gpcOutL0_140);
gpc006 gpcL0_141 ({pp289[5], pp274[3], pp259[1], pp258[5], pp243[3], pp228[1]}, gpcOutL0_141);
gpc006 gpcL0_142 ({pp305[4], pp290[2], pp275[0], pp274[4], pp259[2], pp244[0]}, gpcOutL0_142);
gpc006 gpcL0_143 ({pp305[5], pp290[3], pp275[1], pp274[5], pp259[3], pp244[1]}, gpcOutL0_143);
gpc006 gpcL0_144 ({pp321[4], pp306[2], pp291[0], pp290[4], pp275[2], pp260[0]}, gpcOutL0_144);
gpc006 gpcL0_145 ({pp321[5], pp306[3], pp291[1], pp290[5], pp275[3], pp260[1]}, gpcOutL0_145);
gpc006 gpcL0_146 ({pp337[4], pp322[2], pp307[0], pp306[4], pp291[2], pp276[0]}, gpcOutL0_146);
gpc006 gpcL0_147 ({pp337[5], pp322[3], pp307[1], pp306[5], pp291[3], pp276[1]}, gpcOutL0_147);
gpc006 gpcL0_148 ({pp353[4], pp338[2], pp323[0], pp322[4], pp307[2], pp292[0]}, gpcOutL0_148);
gpc006 gpcL0_149 ({pp353[5], pp338[3], pp323[1], pp322[5], pp307[3], pp292[1]}, gpcOutL0_149);
gpc006 gpcL0_150 ({pp369[4], pp354[2], pp339[0], pp338[4], pp323[2], pp308[0]}, gpcOutL0_150);
gpc006 gpcL0_151 ({pp369[5], pp354[3], pp339[1], pp338[5], pp323[3], pp308[1]}, gpcOutL0_151);
gpc006 gpcL0_152 ({pp385[4], pp370[2], pp355[0], pp354[4], pp339[2], pp324[0]}, gpcOutL0_152);
gpc006 gpcL0_153 ({pp385[5], pp370[3], pp355[1], pp354[5], pp339[3], pp324[1]}, gpcOutL0_153);
gpc006 gpcL0_154 ({pp401[4], pp386[2], pp371[0], pp370[4], pp355[2], pp340[0]}, gpcOutL0_154);
gpc006 gpcL0_155 ({pp401[5], pp386[3], pp371[1], pp370[5], pp355[3], pp340[1]}, gpcOutL0_155);
gpc006 gpcL0_156 ({pp417[4], pp402[2], pp387[0], pp386[4], pp371[2], pp356[0]}, gpcOutL0_156);
gpc006 gpcL0_157 ({pp417[5], pp402[3], pp387[1], pp386[5], pp371[3], pp356[1]}, gpcOutL0_157);
gpc006 gpcL0_158 ({pp433[4], pp418[2], pp403[0], pp402[4], pp387[2], pp372[0]}, gpcOutL0_158);
gpc006 gpcL0_159 ({pp433[5], pp418[3], pp403[1], pp402[5], pp387[3], pp372[1]}, gpcOutL0_159);
gpc006 gpcL0_160 ({pp434[2], pp419[0], pp418[4], pp403[2], pp388[0], pp387[4]}, gpcOutL0_160);
gpc006 gpcL0_161 ({pp434[3], pp419[1], pp418[5], pp403[3], pp388[1], pp387[5]}, gpcOutL0_161);
gpc006 gpcL0_162 ({pp435[0], pp434[4], pp419[2], pp404[0], pp403[4], pp388[2]}, gpcOutL0_162);
gpc006 gpcL0_163 ({pp435[1], pp434[5], pp419[3], pp404[1], pp403[5], pp388[3]}, gpcOutL0_163);
gpc006 gpcL0_164 ({pp435[2], pp420[0], pp419[4], pp404[2], pp389[0], pp388[4]}, gpcOutL0_164);
gpc006 gpcL0_165 ({pp435[3], pp420[1], pp419[5], pp404[3], pp389[1], pp388[5]}, gpcOutL0_165);
gpc006 gpcL0_166 ({pp436[0], pp435[4], pp420[2], pp405[0], pp404[4], pp389[2]}, gpcOutL0_166);
gpc006 gpcL0_167 ({pp436[1], pp435[5], pp420[3], pp405[1], pp404[5], pp389[3]}, gpcOutL0_167);
gpc006 gpcL0_168 ({pp436[2], pp421[0], pp420[4], pp405[2], pp390[0], pp389[4]}, gpcOutL0_168);
gpc006 gpcL0_169 ({pp436[3], pp421[1], pp420[5], pp405[3], pp390[1], pp389[5]}, gpcOutL0_169);
gpc006 gpcL0_170 ({pp437[0], pp436[4], pp421[2], pp406[0], pp405[4], pp390[2]}, gpcOutL0_170);
gpc006 gpcL0_171 ({pp437[1], pp436[5], pp421[3], pp406[1], pp405[5], pp390[3]}, gpcOutL0_171);
gpc006 gpcL0_172 ({pp437[2], pp422[0], pp421[4], pp406[2], pp391[0], pp390[4]}, gpcOutL0_172);
gpc006 gpcL0_173 ({pp437[3], pp422[1], pp421[5], pp406[3], pp391[1], pp390[5]}, gpcOutL0_173);
gpc006 gpcL0_174 ({pp438[0], pp437[4], pp422[2], pp407[0], pp406[4], pp391[2]}, gpcOutL0_174);
gpc006 gpcL0_175 ({pp438[1], pp437[5], pp422[3], pp407[1], pp406[5], pp391[3]}, gpcOutL0_175);
gpc006 gpcL0_176 ({pp438[2], pp423[0], pp422[4], pp407[2], pp392[0], pp391[4]}, gpcOutL0_176);
gpc006 gpcL0_177 ({pp438[3], pp423[1], pp422[5], pp407[3], pp392[1], pp391[5]}, gpcOutL0_177);
gpc006 gpcL0_178 ({pp439[0], pp438[4], pp423[2], pp408[0], pp407[4], pp392[2]}, gpcOutL0_178);
gpc006 gpcL0_179 ({pp439[1], pp438[5], pp423[3], pp408[1], pp407[5], pp392[3]}, gpcOutL0_179);
gpc006 gpcL0_180 ({pp439[2], pp424[0], pp423[4], pp408[2], pp393[0], pp392[4]}, gpcOutL0_180);
gpc006 gpcL0_181 ({pp439[3], pp424[1], pp423[5], pp408[3], pp393[1], pp392[5]}, gpcOutL0_181);
gpc006 gpcL0_182 ({pp440[0], pp439[4], pp424[2], pp409[0], pp408[4], pp393[2]}, gpcOutL0_182);
gpc006 gpcL0_183 ({pp440[1], pp439[5], pp424[3], pp409[1], pp408[5], pp393[3]}, gpcOutL0_183);
gpc006 gpcL0_184 ({pp440[2], pp425[0], pp424[4], pp409[2], pp394[0], pp393[4]}, gpcOutL0_184);
gpc006 gpcL0_185 ({pp440[3], pp425[1], pp424[5], pp409[3], pp394[1], pp393[5]}, gpcOutL0_185);
gpc006 gpcL0_186 ({pp441[0], pp440[4], pp425[2], pp410[0], pp409[4], pp394[2]}, gpcOutL0_186);
gpc006 gpcL0_187 ({pp441[1], pp440[5], pp425[3], pp410[1], pp409[5], pp394[3]}, gpcOutL0_187);
gpc006 gpcL0_188 ({pp441[2], pp426[0], pp425[4], pp410[2], pp395[0], pp394[4]}, gpcOutL0_188);
gpc006 gpcL0_189 ({pp441[3], pp426[1], pp425[5], pp410[3], pp395[1], pp394[5]}, gpcOutL0_189);
gpc006 gpcL0_190 ({pp442[0], pp441[4], pp426[2], pp411[0], pp410[4], pp395[2]}, gpcOutL0_190);
gpc006 gpcL0_191 ({pp442[1], pp441[5], pp426[3], pp411[1], pp410[5], pp395[3]}, gpcOutL0_191);
gpc006 gpcL0_192 ({pp442[2], pp427[0], pp426[4], pp411[2], pp396[0], pp395[4]}, gpcOutL0_192);
gpc006 gpcL0_193 ({pp442[3], pp427[1], pp426[5], pp411[3], pp396[1], pp395[5]}, gpcOutL0_193);
gpc006 gpcL0_194 ({pp443[0], pp442[4], pp427[2], pp412[0], pp411[4], pp396[2]}, gpcOutL0_194);
gpc006 gpcL0_195 ({pp443[1], pp442[5], pp427[3], pp412[1], pp411[5], pp396[3]}, gpcOutL0_195);
gpc006 gpcL0_196 ({pp443[2], pp428[0], pp427[4], pp412[2], pp397[0], pp396[4]}, gpcOutL0_196);
gpc006 gpcL0_197 ({pp443[3], pp428[1], pp427[5], pp412[3], pp397[1], pp396[5]}, gpcOutL0_197);
gpc006 gpcL0_198 ({pp444[0], pp443[4], pp428[2], pp413[0], pp412[4], pp397[2]}, gpcOutL0_198);
gpc006 gpcL0_199 ({pp444[1], pp443[5], pp428[3], pp413[1], pp412[5], pp397[3]}, gpcOutL0_199);
gpc006 gpcL0_200 ({pp444[2], pp429[0], pp428[4], pp413[2], pp398[0], pp397[4]}, gpcOutL0_200);
gpc006 gpcL0_201 ({pp444[3], pp429[1], pp428[5], pp413[3], pp398[1], pp397[5]}, gpcOutL0_201);
gpc006 gpcL0_202 ({pp445[0], pp444[4], pp429[2], pp414[0], pp413[4], pp398[2]}, gpcOutL0_202);
gpc006 gpcL0_203 ({pp445[1], pp444[5], pp429[3], pp414[1], pp413[5], pp398[3]}, gpcOutL0_203);
gpc006 gpcL0_204 ({pp445[2], pp430[0], pp429[4], pp414[2], pp399[0], pp398[4]}, gpcOutL0_204);
gpc006 gpcL0_205 ({pp445[3], pp430[1], pp429[5], pp414[3], pp399[1], pp398[5]}, gpcOutL0_205);
gpc006 gpcL0_206 ({pp446[0], pp445[4], pp430[2], pp415[0], pp414[4], pp399[2]}, gpcOutL0_206);
gpc006 gpcL0_207 ({pp446[1], pp445[5], pp430[3], pp415[1], pp414[5], pp399[3]}, gpcOutL0_207);
gpc006 gpcL0_208 ({pp67[4], pp52[2], pp37[0], pp36[4], pp21[2], pp6[0]}, gpcOutL0_208);
gpc006 gpcL0_209 ({pp67[5], pp52[3], pp37[1], pp36[5], pp21[3], pp6[1]}, gpcOutL0_209);
gpc006 gpcL0_210 ({pp83[4], pp68[2], pp53[0], pp52[4], pp37[2], pp22[0]}, gpcOutL0_210);
gpc006 gpcL0_211 ({pp83[5], pp68[3], pp53[1], pp52[5], pp37[3], pp22[1]}, gpcOutL0_211);
gpc006 gpcL0_212 ({pp99[4], pp84[2], pp69[0], pp68[4], pp53[2], pp38[0]}, gpcOutL0_212);
gpc006 gpcL0_213 ({pp99[5], pp84[3], pp69[1], pp68[5], pp53[3], pp38[1]}, gpcOutL0_213);
gpc006 gpcL0_214 ({pp115[4], pp100[2], pp85[0], pp84[4], pp69[2], pp54[0]}, gpcOutL0_214);
gpc006 gpcL0_215 ({pp115[5], pp100[3], pp85[1], pp84[5], pp69[3], pp54[1]}, gpcOutL0_215);
gpc006 gpcL0_216 ({pp131[4], pp116[2], pp101[0], pp100[4], pp85[2], pp70[0]}, gpcOutL0_216);
gpc006 gpcL0_217 ({pp131[5], pp116[3], pp101[1], pp100[5], pp85[3], pp70[1]}, gpcOutL0_217);
gpc006 gpcL0_218 ({pp147[4], pp132[2], pp117[0], pp116[4], pp101[2], pp86[0]}, gpcOutL0_218);
gpc006 gpcL0_219 ({pp147[5], pp132[3], pp117[1], pp116[5], pp101[3], pp86[1]}, gpcOutL0_219);
gpc006 gpcL0_220 ({pp163[4], pp148[2], pp133[0], pp132[4], pp117[2], pp102[0]}, gpcOutL0_220);
gpc006 gpcL0_221 ({pp163[5], pp148[3], pp133[1], pp132[5], pp117[3], pp102[1]}, gpcOutL0_221);
gpc006 gpcL0_222 ({pp179[4], pp164[2], pp149[0], pp148[4], pp133[2], pp118[0]}, gpcOutL0_222);
gpc006 gpcL0_223 ({pp179[5], pp164[3], pp149[1], pp148[5], pp133[3], pp118[1]}, gpcOutL0_223);
gpc006 gpcL0_224 ({pp195[4], pp180[2], pp165[0], pp164[4], pp149[2], pp134[0]}, gpcOutL0_224);
gpc006 gpcL0_225 ({pp195[5], pp180[3], pp165[1], pp164[5], pp149[3], pp134[1]}, gpcOutL0_225);
gpc006 gpcL0_226 ({pp211[4], pp196[2], pp181[0], pp180[4], pp165[2], pp150[0]}, gpcOutL0_226);
gpc006 gpcL0_227 ({pp211[5], pp196[3], pp181[1], pp180[5], pp165[3], pp150[1]}, gpcOutL0_227);
gpc006 gpcL0_228 ({pp227[4], pp212[2], pp197[0], pp196[4], pp181[2], pp166[0]}, gpcOutL0_228);
gpc006 gpcL0_229 ({pp227[5], pp212[3], pp197[1], pp196[5], pp181[3], pp166[1]}, gpcOutL0_229);
gpc006 gpcL0_230 ({pp243[4], pp228[2], pp213[0], pp212[4], pp197[2], pp182[0]}, gpcOutL0_230);
gpc006 gpcL0_231 ({pp243[5], pp228[3], pp213[1], pp212[5], pp197[3], pp182[1]}, gpcOutL0_231);
gpc006 gpcL0_232 ({pp259[4], pp244[2], pp229[0], pp228[4], pp213[2], pp198[0]}, gpcOutL0_232);
gpc006 gpcL0_233 ({pp259[5], pp244[3], pp229[1], pp228[5], pp213[3], pp198[1]}, gpcOutL0_233);
gpc006 gpcL0_234 ({pp275[4], pp260[2], pp245[0], pp244[4], pp229[2], pp214[0]}, gpcOutL0_234);
gpc006 gpcL0_235 ({pp275[5], pp260[3], pp245[1], pp244[5], pp229[3], pp214[1]}, gpcOutL0_235);
gpc006 gpcL0_236 ({pp291[4], pp276[2], pp261[0], pp260[4], pp245[2], pp230[0]}, gpcOutL0_236);
gpc006 gpcL0_237 ({pp291[5], pp276[3], pp261[1], pp260[5], pp245[3], pp230[1]}, gpcOutL0_237);
gpc006 gpcL0_238 ({pp307[4], pp292[2], pp277[0], pp276[4], pp261[2], pp246[0]}, gpcOutL0_238);
gpc006 gpcL0_239 ({pp307[5], pp292[3], pp277[1], pp276[5], pp261[3], pp246[1]}, gpcOutL0_239);
gpc006 gpcL0_240 ({pp323[4], pp308[2], pp293[0], pp292[4], pp277[2], pp262[0]}, gpcOutL0_240);
gpc006 gpcL0_241 ({pp323[5], pp308[3], pp293[1], pp292[5], pp277[3], pp262[1]}, gpcOutL0_241);
gpc006 gpcL0_242 ({pp339[4], pp324[2], pp309[0], pp308[4], pp293[2], pp278[0]}, gpcOutL0_242);
gpc006 gpcL0_243 ({pp339[5], pp324[3], pp309[1], pp308[5], pp293[3], pp278[1]}, gpcOutL0_243);
gpc006 gpcL0_244 ({pp355[4], pp340[2], pp325[0], pp324[4], pp309[2], pp294[0]}, gpcOutL0_244);
gpc006 gpcL0_245 ({pp355[5], pp340[3], pp325[1], pp324[5], pp309[3], pp294[1]}, gpcOutL0_245);
gpc006 gpcL0_246 ({pp371[4], pp356[2], pp341[0], pp340[4], pp325[2], pp310[0]}, gpcOutL0_246);
gpc006 gpcL0_247 ({pp371[5], pp356[3], pp341[1], pp340[5], pp325[3], pp310[1]}, gpcOutL0_247);
gpc006 gpcL0_248 ({pp372[2], pp357[0], pp356[4], pp341[2], pp326[0], pp325[4]}, gpcOutL0_248);
gpc006 gpcL0_249 ({pp372[3], pp357[1], pp356[5], pp341[3], pp326[1], pp325[5]}, gpcOutL0_249);
gpc006 gpcL0_250 ({pp373[0], pp372[4], pp357[2], pp342[0], pp341[4], pp326[2]}, gpcOutL0_250);
gpc006 gpcL0_251 ({pp373[1], pp372[5], pp357[3], pp342[1], pp341[5], pp326[3]}, gpcOutL0_251);
gpc006 gpcL0_252 ({pp373[2], pp358[0], pp357[4], pp342[2], pp327[0], pp326[4]}, gpcOutL0_252);
gpc006 gpcL0_253 ({pp373[3], pp358[1], pp357[5], pp342[3], pp327[1], pp326[5]}, gpcOutL0_253);
gpc006 gpcL0_254 ({pp374[0], pp373[4], pp358[2], pp343[0], pp342[4], pp327[2]}, gpcOutL0_254);
gpc006 gpcL0_255 ({pp374[1], pp373[5], pp358[3], pp343[1], pp342[5], pp327[3]}, gpcOutL0_255);
gpc006 gpcL0_256 ({pp374[2], pp359[0], pp358[4], pp343[2], pp328[0], pp327[4]}, gpcOutL0_256);
gpc006 gpcL0_257 ({pp374[3], pp359[1], pp358[5], pp343[3], pp328[1], pp327[5]}, gpcOutL0_257);
gpc006 gpcL0_258 ({pp375[0], pp374[4], pp359[2], pp344[0], pp343[4], pp328[2]}, gpcOutL0_258);
gpc006 gpcL0_259 ({pp375[1], pp374[5], pp359[3], pp344[1], pp343[5], pp328[3]}, gpcOutL0_259);
gpc006 gpcL0_260 ({pp375[2], pp360[0], pp359[4], pp344[2], pp329[0], pp328[4]}, gpcOutL0_260);
gpc006 gpcL0_261 ({pp375[3], pp360[1], pp359[5], pp344[3], pp329[1], pp328[5]}, gpcOutL0_261);
gpc006 gpcL0_262 ({pp376[0], pp375[4], pp360[2], pp345[0], pp344[4], pp329[2]}, gpcOutL0_262);
gpc006 gpcL0_263 ({pp376[1], pp375[5], pp360[3], pp345[1], pp344[5], pp329[3]}, gpcOutL0_263);
gpc006 gpcL0_264 ({pp376[2], pp361[0], pp360[4], pp345[2], pp330[0], pp329[4]}, gpcOutL0_264);
gpc006 gpcL0_265 ({pp376[3], pp361[1], pp360[5], pp345[3], pp330[1], pp329[5]}, gpcOutL0_265);
gpc006 gpcL0_266 ({pp377[0], pp376[4], pp361[2], pp346[0], pp345[4], pp330[2]}, gpcOutL0_266);
gpc006 gpcL0_267 ({pp377[1], pp376[5], pp361[3], pp346[1], pp345[5], pp330[3]}, gpcOutL0_267);
gpc006 gpcL0_268 ({pp377[2], pp362[0], pp361[4], pp346[2], pp331[0], pp330[4]}, gpcOutL0_268);
gpc006 gpcL0_269 ({pp377[3], pp362[1], pp361[5], pp346[3], pp331[1], pp330[5]}, gpcOutL0_269);
gpc006 gpcL0_270 ({pp378[0], pp377[4], pp362[2], pp347[0], pp346[4], pp331[2]}, gpcOutL0_270);
gpc006 gpcL0_271 ({pp378[1], pp377[5], pp362[3], pp347[1], pp346[5], pp331[3]}, gpcOutL0_271);
gpc006 gpcL0_272 ({pp378[2], pp363[0], pp362[4], pp347[2], pp332[0], pp331[4]}, gpcOutL0_272);
gpc006 gpcL0_273 ({pp378[3], pp363[1], pp362[5], pp347[3], pp332[1], pp331[5]}, gpcOutL0_273);
gpc006 gpcL0_274 ({pp379[0], pp378[4], pp363[2], pp348[0], pp347[4], pp332[2]}, gpcOutL0_274);
gpc006 gpcL0_275 ({pp379[1], pp378[5], pp363[3], pp348[1], pp347[5], pp332[3]}, gpcOutL0_275);
gpc006 gpcL0_276 ({pp379[2], pp364[0], pp363[4], pp348[2], pp333[0], pp332[4]}, gpcOutL0_276);
gpc006 gpcL0_277 ({pp379[3], pp364[1], pp363[5], pp348[3], pp333[1], pp332[5]}, gpcOutL0_277);
gpc006 gpcL0_278 ({pp380[0], pp379[4], pp364[2], pp349[0], pp348[4], pp333[2]}, gpcOutL0_278);
gpc006 gpcL0_279 ({pp380[1], pp379[5], pp364[3], pp349[1], pp348[5], pp333[3]}, gpcOutL0_279);
gpc006 gpcL0_280 ({pp380[2], pp365[0], pp364[4], pp349[2], pp334[0], pp333[4]}, gpcOutL0_280);
gpc006 gpcL0_281 ({pp380[3], pp365[1], pp364[5], pp349[3], pp334[1], pp333[5]}, gpcOutL0_281);
gpc006 gpcL0_282 ({pp381[0], pp380[4], pp365[2], pp350[0], pp349[4], pp334[2]}, gpcOutL0_282);
gpc006 gpcL0_283 ({pp381[1], pp380[5], pp365[3], pp350[1], pp349[5], pp334[3]}, gpcOutL0_283);
gpc006 gpcL0_284 ({pp381[2], pp366[0], pp365[4], pp350[2], pp335[0], pp334[4]}, gpcOutL0_284);
gpc006 gpcL0_285 ({pp381[3], pp366[1], pp365[5], pp350[3], pp335[1], pp334[5]}, gpcOutL0_285);
gpc006 gpcL0_286 ({pp382[0], pp381[4], pp366[2], pp351[0], pp350[4], pp335[2]}, gpcOutL0_286);
gpc006 gpcL0_287 ({pp382[1], pp381[5], pp366[3], pp351[1], pp350[5], pp335[3]}, gpcOutL0_287);
gpc006 gpcL0_288 ({pp69[4], pp54[2], pp39[0], pp38[4], pp23[2], pp8[0]}, gpcOutL0_288);
gpc006 gpcL0_289 ({pp69[5], pp54[3], pp39[1], pp38[5], pp23[3], pp8[1]}, gpcOutL0_289);
gpc006 gpcL0_290 ({pp85[4], pp70[2], pp55[0], pp54[4], pp39[2], pp24[0]}, gpcOutL0_290);
gpc006 gpcL0_291 ({pp85[5], pp70[3], pp55[1], pp54[5], pp39[3], pp24[1]}, gpcOutL0_291);
gpc006 gpcL0_292 ({pp101[4], pp86[2], pp71[0], pp70[4], pp55[2], pp40[0]}, gpcOutL0_292);
gpc006 gpcL0_293 ({pp101[5], pp86[3], pp71[1], pp70[5], pp55[3], pp40[1]}, gpcOutL0_293);
gpc006 gpcL0_294 ({pp117[4], pp102[2], pp87[0], pp86[4], pp71[2], pp56[0]}, gpcOutL0_294);
gpc006 gpcL0_295 ({pp117[5], pp102[3], pp87[1], pp86[5], pp71[3], pp56[1]}, gpcOutL0_295);
gpc006 gpcL0_296 ({pp133[4], pp118[2], pp103[0], pp102[4], pp87[2], pp72[0]}, gpcOutL0_296);
gpc006 gpcL0_297 ({pp133[5], pp118[3], pp103[1], pp102[5], pp87[3], pp72[1]}, gpcOutL0_297);
gpc006 gpcL0_298 ({pp149[4], pp134[2], pp119[0], pp118[4], pp103[2], pp88[0]}, gpcOutL0_298);
gpc006 gpcL0_299 ({pp149[5], pp134[3], pp119[1], pp118[5], pp103[3], pp88[1]}, gpcOutL0_299);
gpc006 gpcL0_300 ({pp165[4], pp150[2], pp135[0], pp134[4], pp119[2], pp104[0]}, gpcOutL0_300);
gpc006 gpcL0_301 ({pp165[5], pp150[3], pp135[1], pp134[5], pp119[3], pp104[1]}, gpcOutL0_301);
gpc006 gpcL0_302 ({pp181[4], pp166[2], pp151[0], pp150[4], pp135[2], pp120[0]}, gpcOutL0_302);
gpc006 gpcL0_303 ({pp181[5], pp166[3], pp151[1], pp150[5], pp135[3], pp120[1]}, gpcOutL0_303);
gpc006 gpcL0_304 ({pp197[4], pp182[2], pp167[0], pp166[4], pp151[2], pp136[0]}, gpcOutL0_304);
gpc006 gpcL0_305 ({pp197[5], pp182[3], pp167[1], pp166[5], pp151[3], pp136[1]}, gpcOutL0_305);
gpc006 gpcL0_306 ({pp213[4], pp198[2], pp183[0], pp182[4], pp167[2], pp152[0]}, gpcOutL0_306);
gpc006 gpcL0_307 ({pp213[5], pp198[3], pp183[1], pp182[5], pp167[3], pp152[1]}, gpcOutL0_307);
gpc006 gpcL0_308 ({pp229[4], pp214[2], pp199[0], pp198[4], pp183[2], pp168[0]}, gpcOutL0_308);
gpc006 gpcL0_309 ({pp229[5], pp214[3], pp199[1], pp198[5], pp183[3], pp168[1]}, gpcOutL0_309);
gpc006 gpcL0_310 ({pp245[4], pp230[2], pp215[0], pp214[4], pp199[2], pp184[0]}, gpcOutL0_310);
gpc006 gpcL0_311 ({pp245[5], pp230[3], pp215[1], pp214[5], pp199[3], pp184[1]}, gpcOutL0_311);
gpc006 gpcL0_312 ({pp261[4], pp246[2], pp231[0], pp230[4], pp215[2], pp200[0]}, gpcOutL0_312);
gpc006 gpcL0_313 ({pp261[5], pp246[3], pp231[1], pp230[5], pp215[3], pp200[1]}, gpcOutL0_313);
gpc006 gpcL0_314 ({pp277[4], pp262[2], pp247[0], pp246[4], pp231[2], pp216[0]}, gpcOutL0_314);
gpc006 gpcL0_315 ({pp277[5], pp262[3], pp247[1], pp246[5], pp231[3], pp216[1]}, gpcOutL0_315);
gpc006 gpcL0_316 ({pp293[4], pp278[2], pp263[0], pp262[4], pp247[2], pp232[0]}, gpcOutL0_316);
gpc006 gpcL0_317 ({pp293[5], pp278[3], pp263[1], pp262[5], pp247[3], pp232[1]}, gpcOutL0_317);
gpc006 gpcL0_318 ({pp309[4], pp294[2], pp279[0], pp278[4], pp263[2], pp248[0]}, gpcOutL0_318);
gpc006 gpcL0_319 ({pp309[5], pp294[3], pp279[1], pp278[5], pp263[3], pp248[1]}, gpcOutL0_319);
gpc006 gpcL0_320 ({pp310[2], pp295[0], pp294[4], pp279[2], pp264[0], pp263[4]}, gpcOutL0_320);
gpc006 gpcL0_321 ({pp310[3], pp295[1], pp294[5], pp279[3], pp264[1], pp263[5]}, gpcOutL0_321);
gpc006 gpcL0_322 ({pp311[0], pp310[4], pp295[2], pp280[0], pp279[4], pp264[2]}, gpcOutL0_322);
gpc006 gpcL0_323 ({pp311[1], pp310[5], pp295[3], pp280[1], pp279[5], pp264[3]}, gpcOutL0_323);
gpc006 gpcL0_324 ({pp311[2], pp296[0], pp295[4], pp280[2], pp265[0], pp264[4]}, gpcOutL0_324);
gpc006 gpcL0_325 ({pp311[3], pp296[1], pp295[5], pp280[3], pp265[1], pp264[5]}, gpcOutL0_325);
gpc006 gpcL0_326 ({pp312[0], pp311[4], pp296[2], pp281[0], pp280[4], pp265[2]}, gpcOutL0_326);
gpc006 gpcL0_327 ({pp312[1], pp311[5], pp296[3], pp281[1], pp280[5], pp265[3]}, gpcOutL0_327);
gpc006 gpcL0_328 ({pp312[2], pp297[0], pp296[4], pp281[2], pp266[0], pp265[4]}, gpcOutL0_328);
gpc006 gpcL0_329 ({pp312[3], pp297[1], pp296[5], pp281[3], pp266[1], pp265[5]}, gpcOutL0_329);
gpc006 gpcL0_330 ({pp313[0], pp312[4], pp297[2], pp282[0], pp281[4], pp266[2]}, gpcOutL0_330);
gpc006 gpcL0_331 ({pp313[1], pp312[5], pp297[3], pp282[1], pp281[5], pp266[3]}, gpcOutL0_331);
gpc006 gpcL0_332 ({pp313[2], pp298[0], pp297[4], pp282[2], pp267[0], pp266[4]}, gpcOutL0_332);
gpc006 gpcL0_333 ({pp313[3], pp298[1], pp297[5], pp282[3], pp267[1], pp266[5]}, gpcOutL0_333);
gpc006 gpcL0_334 ({pp314[0], pp313[4], pp298[2], pp283[0], pp282[4], pp267[2]}, gpcOutL0_334);
gpc006 gpcL0_335 ({pp314[1], pp313[5], pp298[3], pp283[1], pp282[5], pp267[3]}, gpcOutL0_335);
gpc006 gpcL0_336 ({pp314[2], pp299[0], pp298[4], pp283[2], pp268[0], pp267[4]}, gpcOutL0_336);
gpc006 gpcL0_337 ({pp314[3], pp299[1], pp298[5], pp283[3], pp268[1], pp267[5]}, gpcOutL0_337);
gpc006 gpcL0_338 ({pp315[0], pp314[4], pp299[2], pp284[0], pp283[4], pp268[2]}, gpcOutL0_338);
gpc006 gpcL0_339 ({pp315[1], pp314[5], pp299[3], pp284[1], pp283[5], pp268[3]}, gpcOutL0_339);
gpc006 gpcL0_340 ({pp315[2], pp300[0], pp299[4], pp284[2], pp269[0], pp268[4]}, gpcOutL0_340);
gpc006 gpcL0_341 ({pp315[3], pp300[1], pp299[5], pp284[3], pp269[1], pp268[5]}, gpcOutL0_341);
gpc006 gpcL0_342 ({pp316[0], pp315[4], pp300[2], pp285[0], pp284[4], pp269[2]}, gpcOutL0_342);
gpc006 gpcL0_343 ({pp316[1], pp315[5], pp300[3], pp285[1], pp284[5], pp269[3]}, gpcOutL0_343);
gpc006 gpcL0_344 ({pp316[2], pp301[0], pp300[4], pp285[2], pp270[0], pp269[4]}, gpcOutL0_344);
gpc006 gpcL0_345 ({pp316[3], pp301[1], pp300[5], pp285[3], pp270[1], pp269[5]}, gpcOutL0_345);
gpc006 gpcL0_346 ({pp317[0], pp316[4], pp301[2], pp286[0], pp285[4], pp270[2]}, gpcOutL0_346);
gpc006 gpcL0_347 ({pp317[1], pp316[5], pp301[3], pp286[1], pp285[5], pp270[3]}, gpcOutL0_347);
gpc006 gpcL0_348 ({pp317[2], pp302[0], pp301[4], pp286[2], pp271[0], pp270[4]}, gpcOutL0_348);
gpc006 gpcL0_349 ({pp317[3], pp302[1], pp301[5], pp286[3], pp271[1], pp270[5]}, gpcOutL0_349);
gpc006 gpcL0_350 ({pp318[0], pp317[4], pp302[2], pp287[0], pp286[4], pp271[2]}, gpcOutL0_350);
gpc006 gpcL0_351 ({pp318[1], pp317[5], pp302[3], pp287[1], pp286[5], pp271[3]}, gpcOutL0_351);
gpc006 gpcL0_352 ({pp71[4], pp56[2], pp41[0], pp40[4], pp25[2], pp10[0]}, gpcOutL0_352);
gpc006 gpcL0_353 ({pp71[5], pp56[3], pp41[1], pp40[5], pp25[3], pp10[1]}, gpcOutL0_353);
gpc006 gpcL0_354 ({pp87[4], pp72[2], pp57[0], pp56[4], pp41[2], pp26[0]}, gpcOutL0_354);
gpc006 gpcL0_355 ({pp87[5], pp72[3], pp57[1], pp56[5], pp41[3], pp26[1]}, gpcOutL0_355);
gpc006 gpcL0_356 ({pp103[4], pp88[2], pp73[0], pp72[4], pp57[2], pp42[0]}, gpcOutL0_356);
gpc006 gpcL0_357 ({pp103[5], pp88[3], pp73[1], pp72[5], pp57[3], pp42[1]}, gpcOutL0_357);
gpc006 gpcL0_358 ({pp119[4], pp104[2], pp89[0], pp88[4], pp73[2], pp58[0]}, gpcOutL0_358);
gpc006 gpcL0_359 ({pp119[5], pp104[3], pp89[1], pp88[5], pp73[3], pp58[1]}, gpcOutL0_359);
gpc006 gpcL0_360 ({pp135[4], pp120[2], pp105[0], pp104[4], pp89[2], pp74[0]}, gpcOutL0_360);
gpc006 gpcL0_361 ({pp135[5], pp120[3], pp105[1], pp104[5], pp89[3], pp74[1]}, gpcOutL0_361);
gpc006 gpcL0_362 ({pp151[4], pp136[2], pp121[0], pp120[4], pp105[2], pp90[0]}, gpcOutL0_362);
gpc006 gpcL0_363 ({pp151[5], pp136[3], pp121[1], pp120[5], pp105[3], pp90[1]}, gpcOutL0_363);
gpc006 gpcL0_364 ({pp167[4], pp152[2], pp137[0], pp136[4], pp121[2], pp106[0]}, gpcOutL0_364);
gpc006 gpcL0_365 ({pp167[5], pp152[3], pp137[1], pp136[5], pp121[3], pp106[1]}, gpcOutL0_365);
gpc006 gpcL0_366 ({pp183[4], pp168[2], pp153[0], pp152[4], pp137[2], pp122[0]}, gpcOutL0_366);
gpc006 gpcL0_367 ({pp183[5], pp168[3], pp153[1], pp152[5], pp137[3], pp122[1]}, gpcOutL0_367);
gpc006 gpcL0_368 ({pp199[4], pp184[2], pp169[0], pp168[4], pp153[2], pp138[0]}, gpcOutL0_368);
gpc006 gpcL0_369 ({pp199[5], pp184[3], pp169[1], pp168[5], pp153[3], pp138[1]}, gpcOutL0_369);
gpc006 gpcL0_370 ({pp215[4], pp200[2], pp185[0], pp184[4], pp169[2], pp154[0]}, gpcOutL0_370);
gpc006 gpcL0_371 ({pp215[5], pp200[3], pp185[1], pp184[5], pp169[3], pp154[1]}, gpcOutL0_371);
gpc006 gpcL0_372 ({pp231[4], pp216[2], pp201[0], pp200[4], pp185[2], pp170[0]}, gpcOutL0_372);
gpc006 gpcL0_373 ({pp231[5], pp216[3], pp201[1], pp200[5], pp185[3], pp170[1]}, gpcOutL0_373);
gpc006 gpcL0_374 ({pp247[4], pp232[2], pp217[0], pp216[4], pp201[2], pp186[0]}, gpcOutL0_374);
gpc006 gpcL0_375 ({pp247[5], pp232[3], pp217[1], pp216[5], pp201[3], pp186[1]}, gpcOutL0_375);
gpc006 gpcL0_376 ({pp248[2], pp233[0], pp232[4], pp217[2], pp202[0], pp201[4]}, gpcOutL0_376);
gpc006 gpcL0_377 ({pp248[3], pp233[1], pp232[5], pp217[3], pp202[1], pp201[5]}, gpcOutL0_377);
gpc006 gpcL0_378 ({pp249[0], pp248[4], pp233[2], pp218[0], pp217[4], pp202[2]}, gpcOutL0_378);
gpc006 gpcL0_379 ({pp249[1], pp248[5], pp233[3], pp218[1], pp217[5], pp202[3]}, gpcOutL0_379);
gpc006 gpcL0_380 ({pp249[2], pp234[0], pp233[4], pp218[2], pp203[0], pp202[4]}, gpcOutL0_380);
gpc006 gpcL0_381 ({pp249[3], pp234[1], pp233[5], pp218[3], pp203[1], pp202[5]}, gpcOutL0_381);
gpc006 gpcL0_382 ({pp250[0], pp249[4], pp234[2], pp219[0], pp218[4], pp203[2]}, gpcOutL0_382);
gpc006 gpcL0_383 ({pp250[1], pp249[5], pp234[3], pp219[1], pp218[5], pp203[3]}, gpcOutL0_383);
gpc006 gpcL0_384 ({pp250[2], pp235[0], pp234[4], pp219[2], pp204[0], pp203[4]}, gpcOutL0_384);
gpc006 gpcL0_385 ({pp250[3], pp235[1], pp234[5], pp219[3], pp204[1], pp203[5]}, gpcOutL0_385);
gpc006 gpcL0_386 ({pp251[0], pp250[4], pp235[2], pp220[0], pp219[4], pp204[2]}, gpcOutL0_386);
gpc006 gpcL0_387 ({pp251[1], pp250[5], pp235[3], pp220[1], pp219[5], pp204[3]}, gpcOutL0_387);
gpc006 gpcL0_388 ({pp251[2], pp236[0], pp235[4], pp220[2], pp205[0], pp204[4]}, gpcOutL0_388);
gpc006 gpcL0_389 ({pp251[3], pp236[1], pp235[5], pp220[3], pp205[1], pp204[5]}, gpcOutL0_389);
gpc006 gpcL0_390 ({pp252[0], pp251[4], pp236[2], pp221[0], pp220[4], pp205[2]}, gpcOutL0_390);
gpc006 gpcL0_391 ({pp252[1], pp251[5], pp236[3], pp221[1], pp220[5], pp205[3]}, gpcOutL0_391);
gpc006 gpcL0_392 ({pp252[2], pp237[0], pp236[4], pp221[2], pp206[0], pp205[4]}, gpcOutL0_392);
gpc006 gpcL0_393 ({pp252[3], pp237[1], pp236[5], pp221[3], pp206[1], pp205[5]}, gpcOutL0_393);
gpc006 gpcL0_394 ({pp253[0], pp252[4], pp237[2], pp222[0], pp221[4], pp206[2]}, gpcOutL0_394);
gpc006 gpcL0_395 ({pp253[1], pp252[5], pp237[3], pp222[1], pp221[5], pp206[3]}, gpcOutL0_395);
gpc006 gpcL0_396 ({pp253[2], pp238[0], pp237[4], pp222[2], pp207[0], pp206[4]}, gpcOutL0_396);
gpc006 gpcL0_397 ({pp253[3], pp238[1], pp237[5], pp222[3], pp207[1], pp206[5]}, gpcOutL0_397);
gpc006 gpcL0_398 ({pp254[0], pp253[4], pp238[2], pp223[0], pp222[4], pp207[2]}, gpcOutL0_398);
gpc006 gpcL0_399 ({pp254[1], pp253[5], pp238[3], pp223[1], pp222[5], pp207[3]}, gpcOutL0_399);
gpc006 gpcL0_400 ({pp73[4], pp58[2], pp43[0], pp42[4], pp27[2], pp12[0]}, gpcOutL0_400);
gpc006 gpcL0_401 ({pp73[5], pp58[3], pp43[1], pp42[5], pp27[3], pp12[1]}, gpcOutL0_401);
gpc006 gpcL0_402 ({pp89[4], pp74[2], pp59[0], pp58[4], pp43[2], pp28[0]}, gpcOutL0_402);
gpc006 gpcL0_403 ({pp89[5], pp74[3], pp59[1], pp58[5], pp43[3], pp28[1]}, gpcOutL0_403);
gpc006 gpcL0_404 ({pp105[4], pp90[2], pp75[0], pp74[4], pp59[2], pp44[0]}, gpcOutL0_404);
gpc006 gpcL0_405 ({pp105[5], pp90[3], pp75[1], pp74[5], pp59[3], pp44[1]}, gpcOutL0_405);
gpc006 gpcL0_406 ({pp121[4], pp106[2], pp91[0], pp90[4], pp75[2], pp60[0]}, gpcOutL0_406);
gpc006 gpcL0_407 ({pp121[5], pp106[3], pp91[1], pp90[5], pp75[3], pp60[1]}, gpcOutL0_407);
gpc006 gpcL0_408 ({pp137[4], pp122[2], pp107[0], pp106[4], pp91[2], pp76[0]}, gpcOutL0_408);
gpc006 gpcL0_409 ({pp137[5], pp122[3], pp107[1], pp106[5], pp91[3], pp76[1]}, gpcOutL0_409);
gpc006 gpcL0_410 ({pp153[4], pp138[2], pp123[0], pp122[4], pp107[2], pp92[0]}, gpcOutL0_410);
gpc006 gpcL0_411 ({pp153[5], pp138[3], pp123[1], pp122[5], pp107[3], pp92[1]}, gpcOutL0_411);
gpc006 gpcL0_412 ({pp169[4], pp154[2], pp139[0], pp138[4], pp123[2], pp108[0]}, gpcOutL0_412);
gpc006 gpcL0_413 ({pp169[5], pp154[3], pp139[1], pp138[5], pp123[3], pp108[1]}, gpcOutL0_413);
gpc006 gpcL0_414 ({pp185[4], pp170[2], pp155[0], pp154[4], pp139[2], pp124[0]}, gpcOutL0_414);
gpc006 gpcL0_415 ({pp185[5], pp170[3], pp155[1], pp154[5], pp139[3], pp124[1]}, gpcOutL0_415);
gpc006 gpcL0_416 ({pp186[2], pp171[0], pp170[4], pp155[2], pp140[0], pp139[4]}, gpcOutL0_416);
gpc006 gpcL0_417 ({pp186[3], pp171[1], pp170[5], pp155[3], pp140[1], pp139[5]}, gpcOutL0_417);
gpc006 gpcL0_418 ({pp187[0], pp186[4], pp171[2], pp156[0], pp155[4], pp140[2]}, gpcOutL0_418);
gpc006 gpcL0_419 ({pp187[1], pp186[5], pp171[3], pp156[1], pp155[5], pp140[3]}, gpcOutL0_419);
gpc006 gpcL0_420 ({pp187[2], pp172[0], pp171[4], pp156[2], pp141[0], pp140[4]}, gpcOutL0_420);
gpc006 gpcL0_421 ({pp187[3], pp172[1], pp171[5], pp156[3], pp141[1], pp140[5]}, gpcOutL0_421);
gpc006 gpcL0_422 ({pp188[0], pp187[4], pp172[2], pp157[0], pp156[4], pp141[2]}, gpcOutL0_422);
gpc006 gpcL0_423 ({pp188[1], pp187[5], pp172[3], pp157[1], pp156[5], pp141[3]}, gpcOutL0_423);
gpc006 gpcL0_424 ({pp188[2], pp173[0], pp172[4], pp157[2], pp142[0], pp141[4]}, gpcOutL0_424);
gpc006 gpcL0_425 ({pp188[3], pp173[1], pp172[5], pp157[3], pp142[1], pp141[5]}, gpcOutL0_425);
gpc006 gpcL0_426 ({pp189[0], pp188[4], pp173[2], pp158[0], pp157[4], pp142[2]}, gpcOutL0_426);
gpc006 gpcL0_427 ({pp189[1], pp188[5], pp173[3], pp158[1], pp157[5], pp142[3]}, gpcOutL0_427);
gpc006 gpcL0_428 ({pp189[2], pp174[0], pp173[4], pp158[2], pp143[0], pp142[4]}, gpcOutL0_428);
gpc006 gpcL0_429 ({pp189[3], pp174[1], pp173[5], pp158[3], pp143[1], pp142[5]}, gpcOutL0_429);
gpc006 gpcL0_430 ({pp190[0], pp189[4], pp174[2], pp159[0], pp158[4], pp143[2]}, gpcOutL0_430);
gpc006 gpcL0_431 ({pp190[1], pp189[5], pp174[3], pp159[1], pp158[5], pp143[3]}, gpcOutL0_431);
gpc006 gpcL0_432 ({pp75[4], pp60[2], pp45[0], pp44[4], pp29[2], pp14[0]}, gpcOutL0_432);
gpc006 gpcL0_433 ({pp75[5], pp60[3], pp45[1], pp44[5], pp29[3], pp14[1]}, gpcOutL0_433);
gpc006 gpcL0_434 ({pp91[4], pp76[2], pp61[0], pp60[4], pp45[2], pp30[0]}, gpcOutL0_434);
gpc006 gpcL0_435 ({pp91[5], pp76[3], pp61[1], pp60[5], pp45[3], pp30[1]}, gpcOutL0_435);
gpc006 gpcL0_436 ({pp107[4], pp92[2], pp77[0], pp76[4], pp61[2], pp46[0]}, gpcOutL0_436);
gpc006 gpcL0_437 ({pp107[5], pp92[3], pp77[1], pp76[5], pp61[3], pp46[1]}, gpcOutL0_437);
gpc006 gpcL0_438 ({pp123[4], pp108[2], pp93[0], pp92[4], pp77[2], pp62[0]}, gpcOutL0_438);
gpc006 gpcL0_439 ({pp123[5], pp108[3], pp93[1], pp92[5], pp77[3], pp62[1]}, gpcOutL0_439);
gpc006 gpcL0_440 ({pp124[2], pp109[0], pp108[4], pp93[2], pp78[0], pp77[4]}, gpcOutL0_440);
gpc006 gpcL0_441 ({pp124[3], pp109[1], pp108[5], pp93[3], pp78[1], pp77[5]}, gpcOutL0_441);
gpc006 gpcL0_442 ({pp125[0], pp124[4], pp109[2], pp94[0], pp93[4], pp78[2]}, gpcOutL0_442);
gpc006 gpcL0_443 ({pp125[1], pp124[5], pp109[3], pp94[1], pp93[5], pp78[3]}, gpcOutL0_443);
gpc006 gpcL0_444 ({pp125[2], pp110[0], pp109[4], pp94[2], pp79[0], pp78[4]}, gpcOutL0_444);
gpc006 gpcL0_445 ({pp125[3], pp110[1], pp109[5], pp94[3], pp79[1], pp78[5]}, gpcOutL0_445);
gpc006 gpcL0_446 ({pp126[0], pp125[4], pp110[2], pp95[0], pp94[4], pp79[2]}, gpcOutL0_446);
gpc006 gpcL0_447 ({pp126[1], pp125[5], pp110[3], pp95[1], pp94[5], pp79[3]}, gpcOutL0_447);
gpc015 gpcL0_448 ({pp48[1], pp48[0], pp32[2], pp17[0], pp16[4], pp1[2]}, gpcOutL0_448);
gpc015 gpcL0_449 ({pp49[5], pp49[4], pp34[2], pp19[0], pp18[4], pp3[2]}, gpcOutL0_449);
gpc015 gpcL0_450 ({pp51[5], pp51[4], pp36[2], pp21[0], pp20[4], pp5[2]}, gpcOutL0_450);
gpc015 gpcL0_451 ({pp53[5], pp53[4], pp38[2], pp23[0], pp22[4], pp7[2]}, gpcOutL0_451);
gpc015 gpcL0_452 ({pp55[5], pp55[4], pp40[2], pp25[0], pp24[4], pp9[2]}, gpcOutL0_452);
gpc015 gpcL0_453 ({pp57[5], pp57[4], pp42[2], pp27[0], pp26[4], pp11[2]}, gpcOutL0_453);
gpc015 gpcL0_454 ({pp59[5], pp59[4], pp44[2], pp29[0], pp28[4], pp13[2]}, gpcOutL0_454);
gpc015 gpcL0_455 ({pp61[5], pp61[4], pp46[2], pp31[0], pp30[4], pp15[2]}, gpcOutL0_455);
gpc015 gpcL0_456 ({pp62[3], pp62[2], pp47[0], pp46[4], pp31[2], pp15[4]}, gpcOutL0_456);
gpc015 gpcL0_457 ({pp126[3], pp126[2], pp111[0], pp110[4], pp95[2], pp79[4]}, gpcOutL0_457);
gpc015 gpcL0_458 ({pp190[3], pp190[2], pp175[0], pp174[4], pp159[2], pp143[4]}, gpcOutL0_458);
gpc015 gpcL0_459 ({pp254[3], pp254[2], pp239[0], pp238[4], pp223[2], pp207[4]}, gpcOutL0_459);
gpc015 gpcL0_460 ({pp318[3], pp318[2], pp303[0], pp302[4], pp287[2], pp271[4]}, gpcOutL0_460);
gpc015 gpcL0_461 ({pp382[3], pp382[2], pp367[0], pp366[4], pp351[2], pp335[4]}, gpcOutL0_461);
gpc015 gpcL0_462 ({pp446[3], pp446[2], pp431[0], pp430[4], pp415[2], pp399[4]}, gpcOutL0_462);
gpc015 gpcL0_463 ({pp510[3], pp510[2], pp495[0], pp494[4], pp479[2], pp463[4]}, gpcOutL0_463);
gpc014 gpcL0_464 ({pp32[1], pp32[0], pp16[2], pp1[0], pp0[4]}, gpcOutL0_464);
gpc014 gpcL0_465 ({pp1[4], pp32[3], pp17[1], pp16[5], pp1[3]}, gpcOutL0_465);
gpc014 gpcL0_466 ({pp33[5], pp33[4], pp18[2], pp3[0], pp2[4]}, gpcOutL0_466);
gpc014 gpcL0_467 ({pp3[4], pp34[3], pp19[1], pp18[5], pp3[3]}, gpcOutL0_467);
gpc014 gpcL0_468 ({pp35[5], pp35[4], pp20[2], pp5[0], pp4[4]}, gpcOutL0_468);
gpc014 gpcL0_469 ({pp5[4], pp36[3], pp21[1], pp20[5], pp5[3]}, gpcOutL0_469);
gpc014 gpcL0_470 ({pp37[5], pp37[4], pp22[2], pp7[0], pp6[4]}, gpcOutL0_470);
gpc014 gpcL0_471 ({pp7[4], pp38[3], pp23[1], pp22[5], pp7[3]}, gpcOutL0_471);
gpc014 gpcL0_472 ({pp39[5], pp39[4], pp24[2], pp9[0], pp8[4]}, gpcOutL0_472);
gpc014 gpcL0_473 ({pp9[4], pp40[3], pp25[1], pp24[5], pp9[3]}, gpcOutL0_473);
gpc014 gpcL0_474 ({pp41[5], pp41[4], pp26[2], pp11[0], pp10[4]}, gpcOutL0_474);
gpc014 gpcL0_475 ({pp11[4], pp42[3], pp27[1], pp26[5], pp11[3]}, gpcOutL0_475);
gpc014 gpcL0_476 ({pp43[5], pp43[4], pp28[2], pp13[0], pp12[4]}, gpcOutL0_476);
gpc014 gpcL0_477 ({pp13[4], pp44[3], pp29[1], pp28[5], pp13[3]}, gpcOutL0_477);
gpc014 gpcL0_478 ({pp45[5], pp45[4], pp30[2], pp15[0], pp14[4]}, gpcOutL0_478);
gpc014 gpcL0_479 ({pp63[0], pp47[1], pp46[5], pp31[3], pp15[5]}, gpcOutL0_479);
gpc014 gpcL0_480 ({pp63[2], pp63[1], pp62[5], pp47[3], pp31[5]}, gpcOutL0_480);
gpc014 gpcL0_481 ({pp127[0], pp111[1], pp110[5], pp95[3], pp79[5]}, gpcOutL0_481);
gpc014 gpcL0_482 ({pp127[2], pp127[1], pp126[5], pp111[3], pp95[5]}, gpcOutL0_482);
gpc014 gpcL0_483 ({pp191[0], pp175[1], pp174[5], pp159[3], pp143[5]}, gpcOutL0_483);
gpc014 gpcL0_484 ({pp191[2], pp191[1], pp190[5], pp175[3], pp159[5]}, gpcOutL0_484);
gpc014 gpcL0_485 ({pp255[0], pp239[1], pp238[5], pp223[3], pp207[5]}, gpcOutL0_485);
gpc014 gpcL0_486 ({pp255[2], pp255[1], pp254[5], pp239[3], pp223[5]}, gpcOutL0_486);
gpc014 gpcL0_487 ({pp319[0], pp303[1], pp302[5], pp287[3], pp271[5]}, gpcOutL0_487);
gpc014 gpcL0_488 ({pp319[2], pp319[1], pp318[5], pp303[3], pp287[5]}, gpcOutL0_488);
gpc014 gpcL0_489 ({pp383[0], pp367[1], pp366[5], pp351[3], pp335[5]}, gpcOutL0_489);
gpc014 gpcL0_490 ({pp383[2], pp383[1], pp382[5], pp367[3], pp351[5]}, gpcOutL0_490);
gpc014 gpcL0_491 ({pp447[0], pp431[1], pp430[5], pp415[3], pp399[5]}, gpcOutL0_491);
gpc014 gpcL0_492 ({pp447[2], pp447[1], pp446[5], pp431[3], pp415[5]}, gpcOutL0_492);
gpc014 gpcL0_493 ({pp511[0], pp495[1], pp494[5], pp479[3], pp463[5]}, gpcOutL0_493);
gpc014 gpcL0_494 ({pp511[2], pp511[1], pp510[5], pp495[3], pp479[5]}, gpcOutL0_494);
gpc003 gpcL0_495 ({pp16[3], pp1[1], pp0[5]}, gpcOutL0_495);
gpc003 gpcL0_496 ({pp18[3], pp3[1], pp2[5]}, gpcOutL0_496);
gpc003 gpcL0_497 ({pp20[3], pp5[1], pp4[5]}, gpcOutL0_497);
gpc003 gpcL0_498 ({pp22[3], pp7[1], pp6[5]}, gpcOutL0_498);
gpc003 gpcL0_499 ({pp24[3], pp9[1], pp8[5]}, gpcOutL0_499);
gpc003 gpcL0_500 ({pp26[3], pp11[1], pp10[5]}, gpcOutL0_500);
gpc003 gpcL0_501 ({pp28[3], pp13[1], pp12[5]}, gpcOutL0_501);
gpc003 gpcL0_502 ({pp30[3], pp15[1], pp14[5]}, gpcOutL0_502);
gpc003 gpcL0_503 ({pp46[3], pp31[1], pp30[5]}, gpcOutL0_503);
gpc003 gpcL0_504 ({pp62[4], pp47[2], pp31[4]}, gpcOutL0_504);
gpc003 gpcL0_505 ({pp126[4], pp111[2], pp95[4]}, gpcOutL0_505);
gpc003 gpcL0_506 ({pp190[4], pp175[2], pp159[4]}, gpcOutL0_506);
gpc003 gpcL0_507 ({pp254[4], pp239[2], pp223[4]}, gpcOutL0_507);
gpc003 gpcL0_508 ({pp318[4], pp303[2], pp287[4]}, gpcOutL0_508);
gpc003 gpcL0_509 ({pp382[4], pp367[2], pp351[4]}, gpcOutL0_509);
gpc003 gpcL0_510 ({pp446[4], pp431[2], pp415[4]}, gpcOutL0_510);
gpc003 gpcL0_511 ({pp510[4], pp495[2], pp479[4]}, gpcOutL0_511);
gpc022 gpcL0_512 ({pp17[5], pp2[3], pp17[4], pp2[2]}, gpcOutL0_512);
gpc022 gpcL0_513 ({pp19[5], pp4[3], pp19[4], pp4[2]}, gpcOutL0_513);
gpc022 gpcL0_514 ({pp21[5], pp6[3], pp21[4], pp6[2]}, gpcOutL0_514);
gpc022 gpcL0_515 ({pp23[5], pp8[3], pp23[4], pp8[2]}, gpcOutL0_515);
gpc022 gpcL0_516 ({pp25[5], pp10[3], pp25[4], pp10[2]}, gpcOutL0_516);
gpc022 gpcL0_517 ({pp27[5], pp12[3], pp27[4], pp12[2]}, gpcOutL0_517);
gpc022 gpcL0_518 ({pp29[5], pp14[3], pp29[4], pp14[2]}, gpcOutL0_518);
gpc022 gpcL0_519 ({pp16[1], pp0[3], pp16[0], pp0[2]}, gpcOutL0_519);

// level 1
wire [2:0]  gpcOutL1_0;
wire [2:0]  gpcOutL1_1;
wire [2:0]  gpcOutL1_2;
wire [2:0]  gpcOutL1_3;
wire [2:0]  gpcOutL1_4;
wire [2:0]  gpcOutL1_5;
wire [2:0]  gpcOutL1_6;
wire [2:0]  gpcOutL1_7;
wire [2:0]  gpcOutL1_8;
wire [2:0]  gpcOutL1_9;
wire [2:0]  gpcOutL1_10;
wire [2:0]  gpcOutL1_11;
wire [2:0]  gpcOutL1_12;
wire [2:0]  gpcOutL1_13;
wire [2:0]  gpcOutL1_14;
wire [2:0]  gpcOutL1_15;
wire [2:0]  gpcOutL1_16;
wire [2:0]  gpcOutL1_17;
wire [2:0]  gpcOutL1_18;
wire [2:0]  gpcOutL1_19;
wire [2:0]  gpcOutL1_20;
wire [2:0]  gpcOutL1_21;
wire [2:0]  gpcOutL1_22;
wire [2:0]  gpcOutL1_23;
wire [2:0]  gpcOutL1_24;
wire [2:0]  gpcOutL1_25;
wire [2:0]  gpcOutL1_26;
wire [2:0]  gpcOutL1_27;
wire [2:0]  gpcOutL1_28;
wire [2:0]  gpcOutL1_29;
wire [2:0]  gpcOutL1_30;
wire [2:0]  gpcOutL1_31;
wire [2:0]  gpcOutL1_32;
wire [2:0]  gpcOutL1_33;
wire [2:0]  gpcOutL1_34;
wire [2:0]  gpcOutL1_35;
wire [2:0]  gpcOutL1_36;
wire [2:0]  gpcOutL1_37;
wire [2:0]  gpcOutL1_38;
wire [2:0]  gpcOutL1_39;
wire [2:0]  gpcOutL1_40;
wire [2:0]  gpcOutL1_41;
wire [2:0]  gpcOutL1_42;
wire [2:0]  gpcOutL1_43;
wire [2:0]  gpcOutL1_44;
wire [2:0]  gpcOutL1_45;
wire [2:0]  gpcOutL1_46;
wire [2:0]  gpcOutL1_47;
wire [2:0]  gpcOutL1_48;
wire [2:0]  gpcOutL1_49;
wire [2:0]  gpcOutL1_50;
wire [2:0]  gpcOutL1_51;
wire [2:0]  gpcOutL1_52;
wire [2:0]  gpcOutL1_53;
wire [2:0]  gpcOutL1_54;
wire [2:0]  gpcOutL1_55;
wire [2:0]  gpcOutL1_56;
wire [2:0]  gpcOutL1_57;
wire [2:0]  gpcOutL1_58;
wire [2:0]  gpcOutL1_59;
wire [2:0]  gpcOutL1_60;
wire [2:0]  gpcOutL1_61;
wire [2:0]  gpcOutL1_62;
wire [2:0]  gpcOutL1_63;
wire [2:0]  gpcOutL1_64;
wire [2:0]  gpcOutL1_65;
wire [2:0]  gpcOutL1_66;
wire [2:0]  gpcOutL1_67;
wire [2:0]  gpcOutL1_68;
wire [2:0]  gpcOutL1_69;
wire [2:0]  gpcOutL1_70;
wire [2:0]  gpcOutL1_71;
wire [2:0]  gpcOutL1_72;
wire [2:0]  gpcOutL1_73;
wire [2:0]  gpcOutL1_74;
wire [2:0]  gpcOutL1_75;
wire [2:0]  gpcOutL1_76;
wire [2:0]  gpcOutL1_77;
wire [2:0]  gpcOutL1_78;
wire [2:0]  gpcOutL1_79;
wire [2:0]  gpcOutL1_80;
wire [2:0]  gpcOutL1_81;
wire [2:0]  gpcOutL1_82;
wire [2:0]  gpcOutL1_83;
wire [2:0]  gpcOutL1_84;
wire [2:0]  gpcOutL1_85;
wire [2:0]  gpcOutL1_86;
wire [2:0]  gpcOutL1_87;
wire [2:0]  gpcOutL1_88;
wire [2:0]  gpcOutL1_89;
wire [2:0]  gpcOutL1_90;
wire [2:0]  gpcOutL1_91;
wire [2:0]  gpcOutL1_92;
wire [2:0]  gpcOutL1_93;
wire [2:0]  gpcOutL1_94;
wire [2:0]  gpcOutL1_95;
wire [2:0]  gpcOutL1_96;
wire [2:0]  gpcOutL1_97;
wire [2:0]  gpcOutL1_98;
wire [2:0]  gpcOutL1_99;
wire [2:0]  gpcOutL1_100;
wire [2:0]  gpcOutL1_101;
wire [2:0]  gpcOutL1_102;
wire [2:0]  gpcOutL1_103;
wire [2:0]  gpcOutL1_104;
wire [2:0]  gpcOutL1_105;
wire [2:0]  gpcOutL1_106;
wire [2:0]  gpcOutL1_107;
wire [2:0]  gpcOutL1_108;
wire [2:0]  gpcOutL1_109;
wire [2:0]  gpcOutL1_110;
wire [2:0]  gpcOutL1_111;
wire [2:0]  gpcOutL1_112;
wire [2:0]  gpcOutL1_113;
wire [2:0]  gpcOutL1_114;
wire [2:0]  gpcOutL1_115;
wire [2:0]  gpcOutL1_116;
wire [2:0]  gpcOutL1_117;
wire [2:0]  gpcOutL1_118;
wire [2:0]  gpcOutL1_119;
wire [2:0]  gpcOutL1_120;
wire [2:0]  gpcOutL1_121;
wire [2:0]  gpcOutL1_122;
wire [2:0]  gpcOutL1_123;
wire [2:0]  gpcOutL1_124;
wire [2:0]  gpcOutL1_125;
wire [2:0]  gpcOutL1_126;
wire [2:0]  gpcOutL1_127;
wire [2:0]  gpcOutL1_128;
wire [2:0]  gpcOutL1_129;
wire [2:0]  gpcOutL1_130;
wire [2:0]  gpcOutL1_131;
wire [2:0]  gpcOutL1_132;
wire [2:0]  gpcOutL1_133;
wire [2:0]  gpcOutL1_134;
wire [2:0]  gpcOutL1_135;
wire [2:0]  gpcOutL1_136;
wire [2:0]  gpcOutL1_137;
wire [2:0]  gpcOutL1_138;
wire [2:0]  gpcOutL1_139;
wire [2:0]  gpcOutL1_140;
wire [2:0]  gpcOutL1_141;
wire [2:0]  gpcOutL1_142;
wire [2:0]  gpcOutL1_143;
wire [2:0]  gpcOutL1_144;
wire [2:0]  gpcOutL1_145;
wire [2:0]  gpcOutL1_146;
wire [2:0]  gpcOutL1_147;
wire [2:0]  gpcOutL1_148;
wire [2:0]  gpcOutL1_149;
wire [2:0]  gpcOutL1_150;
wire [2:0]  gpcOutL1_151;
wire [2:0]  gpcOutL1_152;
wire [2:0]  gpcOutL1_153;
wire [2:0]  gpcOutL1_154;
wire [2:0]  gpcOutL1_155;
wire [2:0]  gpcOutL1_156;
wire [2:0]  gpcOutL1_157;
wire [2:0]  gpcOutL1_158;
wire [2:0]  gpcOutL1_159;
wire [2:0]  gpcOutL1_160;
wire [2:0]  gpcOutL1_161;
wire [2:0]  gpcOutL1_162;
wire [2:0]  gpcOutL1_163;
wire [2:0]  gpcOutL1_164;
wire [2:0]  gpcOutL1_165;
wire [2:0]  gpcOutL1_166;
wire [2:0]  gpcOutL1_167;
wire [2:0]  gpcOutL1_168;
wire [2:0]  gpcOutL1_169;
wire [2:0]  gpcOutL1_170;
wire [2:0]  gpcOutL1_171;
wire [2:0]  gpcOutL1_172;
wire [2:0]  gpcOutL1_173;
wire [2:0]  gpcOutL1_174;
wire [2:0]  gpcOutL1_175;
wire [2:0]  gpcOutL1_176;
wire [2:0]  gpcOutL1_177;
wire [2:0]  gpcOutL1_178;
wire [2:0]  gpcOutL1_179;
wire [2:0]  gpcOutL1_180;
wire [2:0]  gpcOutL1_181;
wire [2:0]  gpcOutL1_182;
wire [2:0]  gpcOutL1_183;
wire [2:0]  gpcOutL1_184;
wire [2:0]  gpcOutL1_185;
wire [2:0]  gpcOutL1_186;
wire [2:0]  gpcOutL1_187;
wire [2:0]  gpcOutL1_188;
wire [2:0]  gpcOutL1_189;
wire [2:0]  gpcOutL1_190;
wire [2:0]  gpcOutL1_191;
wire [2:0]  gpcOutL1_192;
wire [2:0]  gpcOutL1_193;
wire [2:0]  gpcOutL1_194;
wire [2:0]  gpcOutL1_195;
wire [2:0]  gpcOutL1_196;
wire [2:0]  gpcOutL1_197;
wire [2:0]  gpcOutL1_198;
wire [2:0]  gpcOutL1_199;
wire [2:0]  gpcOutL1_200;
wire [2:0]  gpcOutL1_201;
wire [2:0]  gpcOutL1_202;
wire [2:0]  gpcOutL1_203;
wire [2:0]  gpcOutL1_204;
wire [2:0]  gpcOutL1_205;
wire [2:0]  gpcOutL1_206;
wire [2:0]  gpcOutL1_207;
wire [2:0]  gpcOutL1_208;
wire [2:0]  gpcOutL1_209;
wire [2:0]  gpcOutL1_210;
wire [2:0]  gpcOutL1_211;
wire [2:0]  gpcOutL1_212;
wire [2:0]  gpcOutL1_213;
wire [2:0]  gpcOutL1_214;
wire [2:0]  gpcOutL1_215;
wire [2:0]  gpcOutL1_216;
wire [2:0]  gpcOutL1_217;
wire [2:0]  gpcOutL1_218;
wire [2:0]  gpcOutL1_219;
wire [2:0]  gpcOutL1_220;
wire [2:0]  gpcOutL1_221;
wire [2:0]  gpcOutL1_222;
wire [2:0]  gpcOutL1_223;
wire [2:0]  gpcOutL1_224;
wire [2:0]  gpcOutL1_225;
wire [2:0]  gpcOutL1_226;
wire [2:0]  gpcOutL1_227;
wire [2:0]  gpcOutL1_228;
wire [2:0]  gpcOutL1_229;
wire [2:0]  gpcOutL1_230;
wire [2:0]  gpcOutL1_231;
wire [2:0]  gpcOutL1_232;
wire [2:0]  gpcOutL1_233;
wire [2:0]  gpcOutL1_234;
wire [2:0]  gpcOutL1_235;
wire [2:0]  gpcOutL1_236;
wire [2:0]  gpcOutL1_237;
wire [2:0]  gpcOutL1_238;
wire [2:0]  gpcOutL1_239;
wire [2:0]  gpcOutL1_240;
wire [2:0]  gpcOutL1_241;
wire [2:0]  gpcOutL1_242;
wire [2:0]  gpcOutL1_243;
wire [2:0]  gpcOutL1_244;
wire [2:0]  gpcOutL1_245;
wire [2:0]  gpcOutL1_246;
wire [2:0]  gpcOutL1_247;
wire [2:0]  gpcOutL1_248;
wire [2:0]  gpcOutL1_249;
wire [2:0]  gpcOutL1_250;
wire [2:0]  gpcOutL1_251;
wire [2:0]  gpcOutL1_252;
wire [2:0]  gpcOutL1_253;
wire [2:0]  gpcOutL1_254;
wire [1:0]  gpcOutL1_255;
wire [1:0]  gpcOutL1_256;
wire [1:0]  gpcOutL1_257;
wire [1:0]  gpcOutL1_258;
wire [1:0]  gpcOutL1_259;
wire [1:0]  gpcOutL1_260;
wire [1:0]  gpcOutL1_261;
wire [1:0]  gpcOutL1_262;
wire [1:0]  gpcOutL1_263;
wire [1:0]  gpcOutL1_264;
wire [1:0]  gpcOutL1_265;
wire [2:0]  gpcOutL1_266;
wire [2:0]  gpcOutL1_267;
wire [2:0]  gpcOutL1_268;
wire [3:0]  gpcOutL1_269;

gpc006 gpcL1_0 ({gpcOutL0_496[1], gpcOutL0_466[2], gpcOutL0_449[0], gpcOutL0_6[0], gpcOutL0_5[1], gpcOutL0_4[2]}, gpcOutL1_0);
gpc006 gpcL1_1 ({gpcOutL0_467[1], gpcOutL0_449[2], gpcOutL0_112[0], gpcOutL0_8[0], gpcOutL0_7[1], gpcOutL0_6[2]}, gpcOutL1_1);
gpc006 gpcL1_2 ({gpcOutL0_467[2], gpcOutL0_113[0], gpcOutL0_112[1], gpcOutL0_9[0], gpcOutL0_8[1], gpcOutL0_7[2]}, gpcOutL1_2);
gpc006 gpcL1_3 ({gpcOutL0_513[0], gpcOutL0_114[0], gpcOutL0_113[1], gpcOutL0_112[2], gpcOutL0_10[0], gpcOutL0_9[1]}, gpcOutL1_3);
gpc006 gpcL1_4 ({gpcOutL0_513[1], gpcOutL0_115[0], gpcOutL0_114[1], gpcOutL0_113[2], gpcOutL0_11[0], gpcOutL0_10[1]}, gpcOutL1_4);
gpc006 gpcL1_5 ({gpcOutL0_513[2], gpcOutL0_468[0], gpcOutL0_116[0], gpcOutL0_115[1], gpcOutL0_114[2], gpcOutL0_12[0]}, gpcOutL1_5);
gpc006 gpcL1_6 ({gpcOutL0_497[0], gpcOutL0_468[1], gpcOutL0_117[0], gpcOutL0_116[1], gpcOutL0_115[2], gpcOutL0_13[0]}, gpcOutL1_6);
gpc006 gpcL1_7 ({gpcOutL0_497[1], gpcOutL0_468[2], gpcOutL0_450[0], gpcOutL0_118[0], gpcOutL0_117[1], gpcOutL0_116[2]}, gpcOutL1_7);
gpc006 gpcL1_8 ({gpcOutL0_469[0], gpcOutL0_450[1], gpcOutL0_119[0], gpcOutL0_118[1], gpcOutL0_117[2], gpcOutL0_15[0]}, gpcOutL1_8);
gpc006 gpcL1_9 ({gpcOutL0_469[1], gpcOutL0_450[2], gpcOutL0_208[0], gpcOutL0_120[0], gpcOutL0_119[1], gpcOutL0_118[2]}, gpcOutL1_9);
gpc006 gpcL1_10 ({gpcOutL0_469[2], gpcOutL0_209[0], gpcOutL0_208[1], gpcOutL0_121[0], gpcOutL0_120[1], gpcOutL0_119[2]}, gpcOutL1_10);
gpc006 gpcL1_11 ({gpcOutL0_514[0], gpcOutL0_210[0], gpcOutL0_209[1], gpcOutL0_208[2], gpcOutL0_122[0], gpcOutL0_121[1]}, gpcOutL1_11);
gpc006 gpcL1_12 ({gpcOutL0_514[1], gpcOutL0_211[0], gpcOutL0_210[1], gpcOutL0_209[2], gpcOutL0_123[0], gpcOutL0_122[1]}, gpcOutL1_12);
gpc006 gpcL1_13 ({gpcOutL0_514[2], gpcOutL0_470[0], gpcOutL0_212[0], gpcOutL0_211[1], gpcOutL0_210[2], gpcOutL0_124[0]}, gpcOutL1_13);
gpc006 gpcL1_14 ({gpcOutL0_498[0], gpcOutL0_470[1], gpcOutL0_213[0], gpcOutL0_212[1], gpcOutL0_211[2], gpcOutL0_125[0]}, gpcOutL1_14);
gpc006 gpcL1_15 ({gpcOutL0_498[1], gpcOutL0_470[2], gpcOutL0_451[0], gpcOutL0_214[0], gpcOutL0_213[1], gpcOutL0_212[2]}, gpcOutL1_15);
gpc006 gpcL1_16 ({gpcOutL0_471[0], gpcOutL0_451[1], gpcOutL0_215[0], gpcOutL0_214[1], gpcOutL0_213[2], gpcOutL0_127[0]}, gpcOutL1_16);
gpc006 gpcL1_17 ({gpcOutL0_471[1], gpcOutL0_451[2], gpcOutL0_288[0], gpcOutL0_216[0], gpcOutL0_215[1], gpcOutL0_214[2]}, gpcOutL1_17);
gpc006 gpcL1_18 ({gpcOutL0_471[2], gpcOutL0_289[0], gpcOutL0_288[1], gpcOutL0_217[0], gpcOutL0_216[1], gpcOutL0_215[2]}, gpcOutL1_18);
gpc006 gpcL1_19 ({gpcOutL0_515[0], gpcOutL0_290[0], gpcOutL0_289[1], gpcOutL0_288[2], gpcOutL0_218[0], gpcOutL0_217[1]}, gpcOutL1_19);
gpc006 gpcL1_20 ({gpcOutL0_515[1], gpcOutL0_291[0], gpcOutL0_290[1], gpcOutL0_289[2], gpcOutL0_219[0], gpcOutL0_218[1]}, gpcOutL1_20);
gpc006 gpcL1_21 ({gpcOutL0_515[2], gpcOutL0_472[0], gpcOutL0_292[0], gpcOutL0_291[1], gpcOutL0_290[2], gpcOutL0_220[0]}, gpcOutL1_21);
gpc006 gpcL1_22 ({gpcOutL0_499[0], gpcOutL0_472[1], gpcOutL0_293[0], gpcOutL0_292[1], gpcOutL0_291[2], gpcOutL0_221[0]}, gpcOutL1_22);
gpc006 gpcL1_23 ({gpcOutL0_499[1], gpcOutL0_472[2], gpcOutL0_452[0], gpcOutL0_294[0], gpcOutL0_293[1], gpcOutL0_292[2]}, gpcOutL1_23);
gpc006 gpcL1_24 ({gpcOutL0_473[0], gpcOutL0_452[1], gpcOutL0_295[0], gpcOutL0_294[1], gpcOutL0_293[2], gpcOutL0_223[0]}, gpcOutL1_24);
gpc006 gpcL1_25 ({gpcOutL0_473[1], gpcOutL0_452[2], gpcOutL0_352[0], gpcOutL0_296[0], gpcOutL0_295[1], gpcOutL0_294[2]}, gpcOutL1_25);
gpc006 gpcL1_26 ({gpcOutL0_473[2], gpcOutL0_353[0], gpcOutL0_352[1], gpcOutL0_297[0], gpcOutL0_296[1], gpcOutL0_295[2]}, gpcOutL1_26);
gpc006 gpcL1_27 ({gpcOutL0_516[0], gpcOutL0_354[0], gpcOutL0_353[1], gpcOutL0_352[2], gpcOutL0_298[0], gpcOutL0_297[1]}, gpcOutL1_27);
gpc006 gpcL1_28 ({gpcOutL0_516[1], gpcOutL0_355[0], gpcOutL0_354[1], gpcOutL0_353[2], gpcOutL0_299[0], gpcOutL0_298[1]}, gpcOutL1_28);
gpc006 gpcL1_29 ({gpcOutL0_516[2], gpcOutL0_474[0], gpcOutL0_356[0], gpcOutL0_355[1], gpcOutL0_354[2], gpcOutL0_300[0]}, gpcOutL1_29);
gpc006 gpcL1_30 ({gpcOutL0_500[0], gpcOutL0_474[1], gpcOutL0_357[0], gpcOutL0_356[1], gpcOutL0_355[2], gpcOutL0_301[0]}, gpcOutL1_30);
gpc006 gpcL1_31 ({gpcOutL0_500[1], gpcOutL0_474[2], gpcOutL0_453[0], gpcOutL0_358[0], gpcOutL0_357[1], gpcOutL0_356[2]}, gpcOutL1_31);
gpc006 gpcL1_32 ({gpcOutL0_475[0], gpcOutL0_453[1], gpcOutL0_359[0], gpcOutL0_358[1], gpcOutL0_357[2], gpcOutL0_303[0]}, gpcOutL1_32);
gpc006 gpcL1_33 ({gpcOutL0_475[1], gpcOutL0_453[2], gpcOutL0_400[0], gpcOutL0_360[0], gpcOutL0_359[1], gpcOutL0_358[2]}, gpcOutL1_33);
gpc006 gpcL1_34 ({gpcOutL0_475[2], gpcOutL0_401[0], gpcOutL0_400[1], gpcOutL0_361[0], gpcOutL0_360[1], gpcOutL0_359[2]}, gpcOutL1_34);
gpc006 gpcL1_35 ({gpcOutL0_517[0], gpcOutL0_402[0], gpcOutL0_401[1], gpcOutL0_400[2], gpcOutL0_362[0], gpcOutL0_361[1]}, gpcOutL1_35);
gpc006 gpcL1_36 ({gpcOutL0_517[1], gpcOutL0_403[0], gpcOutL0_402[1], gpcOutL0_401[2], gpcOutL0_363[0], gpcOutL0_362[1]}, gpcOutL1_36);
gpc006 gpcL1_37 ({gpcOutL0_517[2], gpcOutL0_476[0], gpcOutL0_404[0], gpcOutL0_403[1], gpcOutL0_402[2], gpcOutL0_364[0]}, gpcOutL1_37);
gpc006 gpcL1_38 ({gpcOutL0_501[0], gpcOutL0_476[1], gpcOutL0_405[0], gpcOutL0_404[1], gpcOutL0_403[2], gpcOutL0_365[0]}, gpcOutL1_38);
gpc006 gpcL1_39 ({gpcOutL0_501[1], gpcOutL0_476[2], gpcOutL0_454[0], gpcOutL0_406[0], gpcOutL0_405[1], gpcOutL0_404[2]}, gpcOutL1_39);
gpc006 gpcL1_40 ({gpcOutL0_477[0], gpcOutL0_454[1], gpcOutL0_407[0], gpcOutL0_406[1], gpcOutL0_405[2], gpcOutL0_367[0]}, gpcOutL1_40);
gpc006 gpcL1_41 ({gpcOutL0_477[1], gpcOutL0_454[2], gpcOutL0_432[0], gpcOutL0_408[0], gpcOutL0_407[1], gpcOutL0_406[2]}, gpcOutL1_41);
gpc006 gpcL1_42 ({gpcOutL0_477[2], gpcOutL0_433[0], gpcOutL0_432[1], gpcOutL0_409[0], gpcOutL0_408[1], gpcOutL0_407[2]}, gpcOutL1_42);
gpc006 gpcL1_43 ({gpcOutL0_518[0], gpcOutL0_434[0], gpcOutL0_433[1], gpcOutL0_432[2], gpcOutL0_410[0], gpcOutL0_409[1]}, gpcOutL1_43);
gpc006 gpcL1_44 ({gpcOutL0_518[1], gpcOutL0_435[0], gpcOutL0_434[1], gpcOutL0_433[2], gpcOutL0_411[0], gpcOutL0_410[1]}, gpcOutL1_44);
gpc006 gpcL1_45 ({gpcOutL0_518[2], gpcOutL0_478[0], gpcOutL0_436[0], gpcOutL0_435[1], gpcOutL0_434[2], gpcOutL0_412[0]}, gpcOutL1_45);
gpc006 gpcL1_46 ({gpcOutL0_502[0], gpcOutL0_478[1], gpcOutL0_437[0], gpcOutL0_436[1], gpcOutL0_435[2], gpcOutL0_413[0]}, gpcOutL1_46);
gpc006 gpcL1_47 ({gpcOutL0_502[1], gpcOutL0_478[2], gpcOutL0_455[0], gpcOutL0_438[0], gpcOutL0_437[1], gpcOutL0_436[2]}, gpcOutL1_47);
gpc006 gpcL1_48 ({gpcOutL0_503[0], gpcOutL0_455[1], gpcOutL0_439[0], gpcOutL0_438[1], gpcOutL0_437[2], gpcOutL0_415[0]}, gpcOutL1_48);
gpc006 gpcL1_49 ({gpcOutL0_503[1], gpcOutL0_456[0], gpcOutL0_455[2], gpcOutL0_440[0], gpcOutL0_439[1], gpcOutL0_438[2]}, gpcOutL1_49);
gpc006 gpcL1_50 ({gpcOutL0_479[0], gpcOutL0_456[1], gpcOutL0_441[0], gpcOutL0_440[1], gpcOutL0_439[2], gpcOutL0_417[0]}, gpcOutL1_50);
gpc006 gpcL1_51 ({gpcOutL0_504[0], gpcOutL0_479[1], gpcOutL0_456[2], gpcOutL0_442[0], gpcOutL0_441[1], gpcOutL0_440[2]}, gpcOutL1_51);
gpc006 gpcL1_52 ({gpcOutL0_504[1], gpcOutL0_480[0], gpcOutL0_479[2], gpcOutL0_443[0], gpcOutL0_442[1], gpcOutL0_441[2]}, gpcOutL1_52);
gpc006 gpcL1_53 ({gpcOutL0_480[1], gpcOutL0_444[0], gpcOutL0_443[1], gpcOutL0_442[2], gpcOutL0_420[0], gpcOutL0_419[1]}, gpcOutL1_53);
gpc006 gpcL1_54 ({gpcOutL0_480[2], gpcOutL0_445[0], gpcOutL0_444[1], gpcOutL0_443[2], gpcOutL0_421[0], gpcOutL0_420[1]}, gpcOutL1_54);
gpc006 gpcL1_55 ({gpcOutL0_446[0], gpcOutL0_445[1], gpcOutL0_444[2], gpcOutL0_422[0], gpcOutL0_421[1], gpcOutL0_420[2]}, gpcOutL1_55);
gpc006 gpcL1_56 ({gpcOutL0_447[0], gpcOutL0_446[1], gpcOutL0_445[2], gpcOutL0_423[0], gpcOutL0_422[1], gpcOutL0_421[2]}, gpcOutL1_56);
gpc006 gpcL1_57 ({gpcOutL0_457[0], gpcOutL0_447[1], gpcOutL0_446[2], gpcOutL0_424[0], gpcOutL0_423[1], gpcOutL0_422[2]}, gpcOutL1_57);
gpc006 gpcL1_58 ({gpcOutL0_481[0], gpcOutL0_457[1], gpcOutL0_447[2], gpcOutL0_425[0], gpcOutL0_424[1], gpcOutL0_423[2]}, gpcOutL1_58);
gpc006 gpcL1_59 ({gpcOutL0_505[0], gpcOutL0_481[1], gpcOutL0_457[2], gpcOutL0_426[0], gpcOutL0_425[1], gpcOutL0_424[2]}, gpcOutL1_59);
gpc006 gpcL1_60 ({gpcOutL0_505[1], gpcOutL0_482[0], gpcOutL0_481[2], gpcOutL0_427[0], gpcOutL0_426[1], gpcOutL0_425[2]}, gpcOutL1_60);
gpc006 gpcL1_61 ({gpcOutL0_482[1], gpcOutL0_428[0], gpcOutL0_427[1], gpcOutL0_426[2], gpcOutL0_388[0], gpcOutL0_387[1]}, gpcOutL1_61);
gpc006 gpcL1_62 ({gpcOutL0_482[2], gpcOutL0_429[0], gpcOutL0_428[1], gpcOutL0_427[2], gpcOutL0_389[0], gpcOutL0_388[1]}, gpcOutL1_62);
gpc006 gpcL1_63 ({gpcOutL0_430[0], gpcOutL0_429[1], gpcOutL0_428[2], gpcOutL0_390[0], gpcOutL0_389[1], gpcOutL0_388[2]}, gpcOutL1_63);
gpc006 gpcL1_64 ({gpcOutL0_431[0], gpcOutL0_430[1], gpcOutL0_429[2], gpcOutL0_391[0], gpcOutL0_390[1], gpcOutL0_389[2]}, gpcOutL1_64);
gpc006 gpcL1_65 ({gpcOutL0_458[0], gpcOutL0_431[1], gpcOutL0_430[2], gpcOutL0_392[0], gpcOutL0_391[1], gpcOutL0_390[2]}, gpcOutL1_65);
gpc006 gpcL1_66 ({gpcOutL0_483[0], gpcOutL0_458[1], gpcOutL0_431[2], gpcOutL0_393[0], gpcOutL0_392[1], gpcOutL0_391[2]}, gpcOutL1_66);
gpc006 gpcL1_67 ({gpcOutL0_506[0], gpcOutL0_483[1], gpcOutL0_458[2], gpcOutL0_394[0], gpcOutL0_393[1], gpcOutL0_392[2]}, gpcOutL1_67);
gpc006 gpcL1_68 ({gpcOutL0_506[1], gpcOutL0_484[0], gpcOutL0_483[2], gpcOutL0_395[0], gpcOutL0_394[1], gpcOutL0_393[2]}, gpcOutL1_68);
gpc006 gpcL1_69 ({gpcOutL0_484[1], gpcOutL0_396[0], gpcOutL0_395[1], gpcOutL0_394[2], gpcOutL0_340[0], gpcOutL0_339[1]}, gpcOutL1_69);
gpc006 gpcL1_70 ({gpcOutL0_484[2], gpcOutL0_397[0], gpcOutL0_396[1], gpcOutL0_395[2], gpcOutL0_341[0], gpcOutL0_340[1]}, gpcOutL1_70);
gpc006 gpcL1_71 ({gpcOutL0_398[0], gpcOutL0_397[1], gpcOutL0_396[2], gpcOutL0_342[0], gpcOutL0_341[1], gpcOutL0_340[2]}, gpcOutL1_71);
gpc006 gpcL1_72 ({gpcOutL0_399[0], gpcOutL0_398[1], gpcOutL0_397[2], gpcOutL0_343[0], gpcOutL0_342[1], gpcOutL0_341[2]}, gpcOutL1_72);
gpc006 gpcL1_73 ({gpcOutL0_459[0], gpcOutL0_399[1], gpcOutL0_398[2], gpcOutL0_344[0], gpcOutL0_343[1], gpcOutL0_342[2]}, gpcOutL1_73);
gpc006 gpcL1_74 ({gpcOutL0_485[0], gpcOutL0_459[1], gpcOutL0_399[2], gpcOutL0_345[0], gpcOutL0_344[1], gpcOutL0_343[2]}, gpcOutL1_74);
gpc006 gpcL1_75 ({gpcOutL0_507[0], gpcOutL0_485[1], gpcOutL0_459[2], gpcOutL0_346[0], gpcOutL0_345[1], gpcOutL0_344[2]}, gpcOutL1_75);
gpc006 gpcL1_76 ({gpcOutL0_507[1], gpcOutL0_486[0], gpcOutL0_485[2], gpcOutL0_347[0], gpcOutL0_346[1], gpcOutL0_345[2]}, gpcOutL1_76);
gpc006 gpcL1_77 ({gpcOutL0_486[1], gpcOutL0_348[0], gpcOutL0_347[1], gpcOutL0_346[2], gpcOutL0_276[0], gpcOutL0_275[1]}, gpcOutL1_77);
gpc006 gpcL1_78 ({gpcOutL0_486[2], gpcOutL0_349[0], gpcOutL0_348[1], gpcOutL0_347[2], gpcOutL0_277[0], gpcOutL0_276[1]}, gpcOutL1_78);
gpc006 gpcL1_79 ({gpcOutL0_350[0], gpcOutL0_349[1], gpcOutL0_348[2], gpcOutL0_278[0], gpcOutL0_277[1], gpcOutL0_276[2]}, gpcOutL1_79);
gpc006 gpcL1_80 ({gpcOutL0_351[0], gpcOutL0_350[1], gpcOutL0_349[2], gpcOutL0_279[0], gpcOutL0_278[1], gpcOutL0_277[2]}, gpcOutL1_80);
gpc006 gpcL1_81 ({gpcOutL0_460[0], gpcOutL0_351[1], gpcOutL0_350[2], gpcOutL0_280[0], gpcOutL0_279[1], gpcOutL0_278[2]}, gpcOutL1_81);
gpc006 gpcL1_82 ({gpcOutL0_487[0], gpcOutL0_460[1], gpcOutL0_351[2], gpcOutL0_281[0], gpcOutL0_280[1], gpcOutL0_279[2]}, gpcOutL1_82);
gpc006 gpcL1_83 ({gpcOutL0_508[0], gpcOutL0_487[1], gpcOutL0_460[2], gpcOutL0_282[0], gpcOutL0_281[1], gpcOutL0_280[2]}, gpcOutL1_83);
gpc006 gpcL1_84 ({gpcOutL0_508[1], gpcOutL0_488[0], gpcOutL0_487[2], gpcOutL0_283[0], gpcOutL0_282[1], gpcOutL0_281[2]}, gpcOutL1_84);
gpc006 gpcL1_85 ({gpcOutL0_488[1], gpcOutL0_284[0], gpcOutL0_283[1], gpcOutL0_282[2], gpcOutL0_196[0], gpcOutL0_195[1]}, gpcOutL1_85);
gpc006 gpcL1_86 ({gpcOutL0_488[2], gpcOutL0_285[0], gpcOutL0_284[1], gpcOutL0_283[2], gpcOutL0_197[0], gpcOutL0_196[1]}, gpcOutL1_86);
gpc006 gpcL1_87 ({gpcOutL0_286[0], gpcOutL0_285[1], gpcOutL0_284[2], gpcOutL0_198[0], gpcOutL0_197[1], gpcOutL0_196[2]}, gpcOutL1_87);
gpc006 gpcL1_88 ({gpcOutL0_287[0], gpcOutL0_286[1], gpcOutL0_285[2], gpcOutL0_199[0], gpcOutL0_198[1], gpcOutL0_197[2]}, gpcOutL1_88);
gpc006 gpcL1_89 ({gpcOutL0_461[0], gpcOutL0_287[1], gpcOutL0_286[2], gpcOutL0_200[0], gpcOutL0_199[1], gpcOutL0_198[2]}, gpcOutL1_89);
gpc006 gpcL1_90 ({gpcOutL0_489[0], gpcOutL0_461[1], gpcOutL0_287[2], gpcOutL0_201[0], gpcOutL0_200[1], gpcOutL0_199[2]}, gpcOutL1_90);
gpc006 gpcL1_91 ({gpcOutL0_509[0], gpcOutL0_489[1], gpcOutL0_461[2], gpcOutL0_202[0], gpcOutL0_201[1], gpcOutL0_200[2]}, gpcOutL1_91);
gpc006 gpcL1_92 ({gpcOutL0_509[1], gpcOutL0_490[0], gpcOutL0_489[2], gpcOutL0_203[0], gpcOutL0_202[1], gpcOutL0_201[2]}, gpcOutL1_92);
gpc006 gpcL1_93 ({gpcOutL0_490[1], gpcOutL0_204[0], gpcOutL0_203[1], gpcOutL0_202[2], gpcOutL0_100[0], gpcOutL0_99[1]}, gpcOutL1_93);
gpc006 gpcL1_94 ({gpcOutL0_490[2], gpcOutL0_205[0], gpcOutL0_204[1], gpcOutL0_203[2], gpcOutL0_101[0], gpcOutL0_100[1]}, gpcOutL1_94);
gpc006 gpcL1_95 ({gpcOutL0_206[0], gpcOutL0_205[1], gpcOutL0_204[2], gpcOutL0_102[0], gpcOutL0_101[1], gpcOutL0_100[2]}, gpcOutL1_95);
gpc006 gpcL1_96 ({gpcOutL0_207[0], gpcOutL0_206[1], gpcOutL0_205[2], gpcOutL0_103[0], gpcOutL0_102[1], gpcOutL0_101[2]}, gpcOutL1_96);
gpc006 gpcL1_97 ({gpcOutL0_462[0], gpcOutL0_207[1], gpcOutL0_206[2], gpcOutL0_104[0], gpcOutL0_103[1], gpcOutL0_102[2]}, gpcOutL1_97);
gpc006 gpcL1_98 ({gpcOutL0_491[0], gpcOutL0_462[1], gpcOutL0_207[2], gpcOutL0_105[0], gpcOutL0_104[1], gpcOutL0_103[2]}, gpcOutL1_98);
gpc006 gpcL1_99 ({gpcOutL0_510[0], gpcOutL0_491[1], gpcOutL0_462[2], gpcOutL0_106[0], gpcOutL0_105[1], gpcOutL0_104[2]}, gpcOutL1_99);
gpc006 gpcL1_100 ({gpcOutL0_510[1], gpcOutL0_492[0], gpcOutL0_491[2], gpcOutL0_107[0], gpcOutL0_106[1], gpcOutL0_105[2]}, gpcOutL1_100);
gpc006 gpcL1_101 ({gpcOutL0_492[2], gpcOutL0_109[0], gpcOutL0_108[1], gpcOutL0_107[2], pp447[3], pp431[5]}, gpcOutL1_101);
gpc006 gpcL1_102 ({gpcOutL0_126[0], gpcOutL0_125[1], gpcOutL0_124[2], gpcOutL0_22[0], gpcOutL0_21[1], gpcOutL0_20[2]}, gpcOutL1_102);
gpc006 gpcL1_103 ({gpcOutL0_128[0], gpcOutL0_127[1], gpcOutL0_126[2], gpcOutL0_24[0], gpcOutL0_23[1], gpcOutL0_22[2]}, gpcOutL1_103);
gpc006 gpcL1_104 ({gpcOutL0_129[0], gpcOutL0_128[1], gpcOutL0_127[2], gpcOutL0_25[0], gpcOutL0_24[1], gpcOutL0_23[2]}, gpcOutL1_104);
gpc006 gpcL1_105 ({gpcOutL0_216[2], gpcOutL0_130[0], gpcOutL0_129[1], gpcOutL0_128[2], gpcOutL0_26[0], gpcOutL0_25[1]}, gpcOutL1_105);
gpc006 gpcL1_106 ({gpcOutL0_217[2], gpcOutL0_131[0], gpcOutL0_130[1], gpcOutL0_129[2], gpcOutL0_27[0], gpcOutL0_26[1]}, gpcOutL1_106);
gpc006 gpcL1_107 ({gpcOutL0_219[1], gpcOutL0_218[2], gpcOutL0_132[0], gpcOutL0_131[1], gpcOutL0_130[2], gpcOutL0_28[0]}, gpcOutL1_107);
gpc006 gpcL1_108 ({gpcOutL0_220[1], gpcOutL0_219[2], gpcOutL0_133[0], gpcOutL0_132[1], gpcOutL0_131[2], gpcOutL0_29[0]}, gpcOutL1_108);
gpc006 gpcL1_109 ({gpcOutL0_222[0], gpcOutL0_221[1], gpcOutL0_220[2], gpcOutL0_134[0], gpcOutL0_133[1], gpcOutL0_132[2]}, gpcOutL1_109);
gpc006 gpcL1_110 ({gpcOutL0_222[1], gpcOutL0_221[2], gpcOutL0_135[0], gpcOutL0_134[1], gpcOutL0_133[2], gpcOutL0_31[0]}, gpcOutL1_110);
gpc006 gpcL1_111 ({gpcOutL0_224[0], gpcOutL0_223[1], gpcOutL0_222[2], gpcOutL0_136[0], gpcOutL0_135[1], gpcOutL0_134[2]}, gpcOutL1_111);
gpc006 gpcL1_112 ({gpcOutL0_225[0], gpcOutL0_224[1], gpcOutL0_223[2], gpcOutL0_137[0], gpcOutL0_136[1], gpcOutL0_135[2]}, gpcOutL1_112);
gpc006 gpcL1_113 ({gpcOutL0_296[2], gpcOutL0_226[0], gpcOutL0_225[1], gpcOutL0_224[2], gpcOutL0_138[0], gpcOutL0_137[1]}, gpcOutL1_113);
gpc006 gpcL1_114 ({gpcOutL0_297[2], gpcOutL0_227[0], gpcOutL0_226[1], gpcOutL0_225[2], gpcOutL0_139[0], gpcOutL0_138[1]}, gpcOutL1_114);
gpc006 gpcL1_115 ({gpcOutL0_299[1], gpcOutL0_298[2], gpcOutL0_228[0], gpcOutL0_227[1], gpcOutL0_226[2], gpcOutL0_140[0]}, gpcOutL1_115);
gpc006 gpcL1_116 ({gpcOutL0_300[1], gpcOutL0_299[2], gpcOutL0_229[0], gpcOutL0_228[1], gpcOutL0_227[2], gpcOutL0_141[0]}, gpcOutL1_116);
gpc006 gpcL1_117 ({gpcOutL0_302[0], gpcOutL0_301[1], gpcOutL0_300[2], gpcOutL0_230[0], gpcOutL0_229[1], gpcOutL0_228[2]}, gpcOutL1_117);
gpc006 gpcL1_118 ({gpcOutL0_302[1], gpcOutL0_301[2], gpcOutL0_231[0], gpcOutL0_230[1], gpcOutL0_229[2], gpcOutL0_143[0]}, gpcOutL1_118);
gpc006 gpcL1_119 ({gpcOutL0_304[0], gpcOutL0_303[1], gpcOutL0_302[2], gpcOutL0_232[0], gpcOutL0_231[1], gpcOutL0_230[2]}, gpcOutL1_119);
gpc006 gpcL1_120 ({gpcOutL0_305[0], gpcOutL0_304[1], gpcOutL0_303[2], gpcOutL0_233[0], gpcOutL0_232[1], gpcOutL0_231[2]}, gpcOutL1_120);
gpc006 gpcL1_121 ({gpcOutL0_360[2], gpcOutL0_306[0], gpcOutL0_305[1], gpcOutL0_304[2], gpcOutL0_234[0], gpcOutL0_233[1]}, gpcOutL1_121);
gpc006 gpcL1_122 ({gpcOutL0_361[2], gpcOutL0_307[0], gpcOutL0_306[1], gpcOutL0_305[2], gpcOutL0_235[0], gpcOutL0_234[1]}, gpcOutL1_122);
gpc006 gpcL1_123 ({gpcOutL0_363[1], gpcOutL0_362[2], gpcOutL0_308[0], gpcOutL0_307[1], gpcOutL0_306[2], gpcOutL0_236[0]}, gpcOutL1_123);
gpc006 gpcL1_124 ({gpcOutL0_364[1], gpcOutL0_363[2], gpcOutL0_309[0], gpcOutL0_308[1], gpcOutL0_307[2], gpcOutL0_237[0]}, gpcOutL1_124);
gpc006 gpcL1_125 ({gpcOutL0_366[0], gpcOutL0_365[1], gpcOutL0_364[2], gpcOutL0_310[0], gpcOutL0_309[1], gpcOutL0_308[2]}, gpcOutL1_125);
gpc006 gpcL1_126 ({gpcOutL0_366[1], gpcOutL0_365[2], gpcOutL0_311[0], gpcOutL0_310[1], gpcOutL0_309[2], gpcOutL0_239[0]}, gpcOutL1_126);
gpc006 gpcL1_127 ({gpcOutL0_368[0], gpcOutL0_367[1], gpcOutL0_366[2], gpcOutL0_312[0], gpcOutL0_311[1], gpcOutL0_310[2]}, gpcOutL1_127);
gpc006 gpcL1_128 ({gpcOutL0_369[0], gpcOutL0_368[1], gpcOutL0_367[2], gpcOutL0_313[0], gpcOutL0_312[1], gpcOutL0_311[2]}, gpcOutL1_128);
gpc006 gpcL1_129 ({gpcOutL0_408[2], gpcOutL0_370[0], gpcOutL0_369[1], gpcOutL0_368[2], gpcOutL0_314[0], gpcOutL0_313[1]}, gpcOutL1_129);
gpc006 gpcL1_130 ({gpcOutL0_409[2], gpcOutL0_371[0], gpcOutL0_370[1], gpcOutL0_369[2], gpcOutL0_315[0], gpcOutL0_314[1]}, gpcOutL1_130);
gpc006 gpcL1_131 ({gpcOutL0_411[1], gpcOutL0_410[2], gpcOutL0_372[0], gpcOutL0_371[1], gpcOutL0_370[2], gpcOutL0_316[0]}, gpcOutL1_131);
gpc006 gpcL1_132 ({gpcOutL0_412[1], gpcOutL0_411[2], gpcOutL0_373[0], gpcOutL0_372[1], gpcOutL0_371[2], gpcOutL0_317[0]}, gpcOutL1_132);
gpc006 gpcL1_133 ({gpcOutL0_414[0], gpcOutL0_413[1], gpcOutL0_412[2], gpcOutL0_374[0], gpcOutL0_373[1], gpcOutL0_372[2]}, gpcOutL1_133);
gpc006 gpcL1_134 ({gpcOutL0_414[1], gpcOutL0_413[2], gpcOutL0_375[0], gpcOutL0_374[1], gpcOutL0_373[2], gpcOutL0_319[0]}, gpcOutL1_134);
gpc006 gpcL1_135 ({gpcOutL0_416[0], gpcOutL0_415[1], gpcOutL0_414[2], gpcOutL0_376[0], gpcOutL0_375[1], gpcOutL0_374[2]}, gpcOutL1_135);
gpc006 gpcL1_136 ({gpcOutL0_416[1], gpcOutL0_415[2], gpcOutL0_377[0], gpcOutL0_376[1], gpcOutL0_375[2], gpcOutL0_321[0]}, gpcOutL1_136);
gpc006 gpcL1_137 ({gpcOutL0_418[0], gpcOutL0_417[1], gpcOutL0_416[2], gpcOutL0_378[0], gpcOutL0_377[1], gpcOutL0_376[2]}, gpcOutL1_137);
gpc006 gpcL1_138 ({gpcOutL0_419[0], gpcOutL0_418[1], gpcOutL0_417[2], gpcOutL0_379[0], gpcOutL0_378[1], gpcOutL0_377[2]}, gpcOutL1_138);
gpc006 gpcL1_139 ({gpcOutL0_418[2], gpcOutL0_380[0], gpcOutL0_379[1], gpcOutL0_378[2], gpcOutL0_324[0], gpcOutL0_323[1]}, gpcOutL1_139);
gpc006 gpcL1_140 ({gpcOutL0_419[2], gpcOutL0_381[0], gpcOutL0_380[1], gpcOutL0_379[2], gpcOutL0_325[0], gpcOutL0_324[1]}, gpcOutL1_140);
gpc006 gpcL1_141 ({gpcOutL0_382[0], gpcOutL0_381[1], gpcOutL0_380[2], gpcOutL0_326[0], gpcOutL0_325[1], gpcOutL0_324[2]}, gpcOutL1_141);
gpc006 gpcL1_142 ({gpcOutL0_383[0], gpcOutL0_382[1], gpcOutL0_381[2], gpcOutL0_327[0], gpcOutL0_326[1], gpcOutL0_325[2]}, gpcOutL1_142);
gpc006 gpcL1_143 ({gpcOutL0_384[0], gpcOutL0_383[1], gpcOutL0_382[2], gpcOutL0_328[0], gpcOutL0_327[1], gpcOutL0_326[2]}, gpcOutL1_143);
gpc006 gpcL1_144 ({gpcOutL0_385[0], gpcOutL0_384[1], gpcOutL0_383[2], gpcOutL0_329[0], gpcOutL0_328[1], gpcOutL0_327[2]}, gpcOutL1_144);
gpc006 gpcL1_145 ({gpcOutL0_386[0], gpcOutL0_385[1], gpcOutL0_384[2], gpcOutL0_330[0], gpcOutL0_329[1], gpcOutL0_328[2]}, gpcOutL1_145);
gpc006 gpcL1_146 ({gpcOutL0_387[0], gpcOutL0_386[1], gpcOutL0_385[2], gpcOutL0_331[0], gpcOutL0_330[1], gpcOutL0_329[2]}, gpcOutL1_146);
gpc006 gpcL1_147 ({gpcOutL0_386[2], gpcOutL0_332[0], gpcOutL0_331[1], gpcOutL0_330[2], gpcOutL0_260[0], gpcOutL0_259[1]}, gpcOutL1_147);
gpc006 gpcL1_148 ({gpcOutL0_387[2], gpcOutL0_333[0], gpcOutL0_332[1], gpcOutL0_331[2], gpcOutL0_261[0], gpcOutL0_260[1]}, gpcOutL1_148);
gpc006 gpcL1_149 ({gpcOutL0_334[0], gpcOutL0_333[1], gpcOutL0_332[2], gpcOutL0_262[0], gpcOutL0_261[1], gpcOutL0_260[2]}, gpcOutL1_149);
gpc006 gpcL1_150 ({gpcOutL0_335[0], gpcOutL0_334[1], gpcOutL0_333[2], gpcOutL0_263[0], gpcOutL0_262[1], gpcOutL0_261[2]}, gpcOutL1_150);
gpc006 gpcL1_151 ({gpcOutL0_336[0], gpcOutL0_335[1], gpcOutL0_334[2], gpcOutL0_264[0], gpcOutL0_263[1], gpcOutL0_262[2]}, gpcOutL1_151);
gpc006 gpcL1_152 ({gpcOutL0_337[0], gpcOutL0_336[1], gpcOutL0_335[2], gpcOutL0_265[0], gpcOutL0_264[1], gpcOutL0_263[2]}, gpcOutL1_152);
gpc006 gpcL1_153 ({gpcOutL0_338[0], gpcOutL0_337[1], gpcOutL0_336[2], gpcOutL0_266[0], gpcOutL0_265[1], gpcOutL0_264[2]}, gpcOutL1_153);
gpc006 gpcL1_154 ({gpcOutL0_339[0], gpcOutL0_338[1], gpcOutL0_337[2], gpcOutL0_267[0], gpcOutL0_266[1], gpcOutL0_265[2]}, gpcOutL1_154);
gpc006 gpcL1_155 ({gpcOutL0_338[2], gpcOutL0_268[0], gpcOutL0_267[1], gpcOutL0_266[2], gpcOutL0_180[0], gpcOutL0_179[1]}, gpcOutL1_155);
gpc006 gpcL1_156 ({gpcOutL0_339[2], gpcOutL0_269[0], gpcOutL0_268[1], gpcOutL0_267[2], gpcOutL0_181[0], gpcOutL0_180[1]}, gpcOutL1_156);
gpc006 gpcL1_157 ({gpcOutL0_270[0], gpcOutL0_269[1], gpcOutL0_268[2], gpcOutL0_182[0], gpcOutL0_181[1], gpcOutL0_180[2]}, gpcOutL1_157);
gpc006 gpcL1_158 ({gpcOutL0_271[0], gpcOutL0_270[1], gpcOutL0_269[2], gpcOutL0_183[0], gpcOutL0_182[1], gpcOutL0_181[2]}, gpcOutL1_158);
gpc006 gpcL1_159 ({gpcOutL0_272[0], gpcOutL0_271[1], gpcOutL0_270[2], gpcOutL0_184[0], gpcOutL0_183[1], gpcOutL0_182[2]}, gpcOutL1_159);
gpc006 gpcL1_160 ({gpcOutL0_273[0], gpcOutL0_272[1], gpcOutL0_271[2], gpcOutL0_185[0], gpcOutL0_184[1], gpcOutL0_183[2]}, gpcOutL1_160);
gpc006 gpcL1_161 ({gpcOutL0_274[0], gpcOutL0_273[1], gpcOutL0_272[2], gpcOutL0_186[0], gpcOutL0_185[1], gpcOutL0_184[2]}, gpcOutL1_161);
gpc006 gpcL1_162 ({gpcOutL0_275[0], gpcOutL0_274[1], gpcOutL0_273[2], gpcOutL0_187[0], gpcOutL0_186[1], gpcOutL0_185[2]}, gpcOutL1_162);
gpc006 gpcL1_163 ({gpcOutL0_274[2], gpcOutL0_188[0], gpcOutL0_187[1], gpcOutL0_186[2], gpcOutL0_84[0], gpcOutL0_83[1]}, gpcOutL1_163);
gpc006 gpcL1_164 ({gpcOutL0_275[2], gpcOutL0_189[0], gpcOutL0_188[1], gpcOutL0_187[2], gpcOutL0_85[0], gpcOutL0_84[1]}, gpcOutL1_164);
gpc006 gpcL1_165 ({gpcOutL0_190[0], gpcOutL0_189[1], gpcOutL0_188[2], gpcOutL0_86[0], gpcOutL0_85[1], gpcOutL0_84[2]}, gpcOutL1_165);
gpc006 gpcL1_166 ({gpcOutL0_191[0], gpcOutL0_190[1], gpcOutL0_189[2], gpcOutL0_87[0], gpcOutL0_86[1], gpcOutL0_85[2]}, gpcOutL1_166);
gpc006 gpcL1_167 ({gpcOutL0_192[0], gpcOutL0_191[1], gpcOutL0_190[2], gpcOutL0_88[0], gpcOutL0_87[1], gpcOutL0_86[2]}, gpcOutL1_167);
gpc006 gpcL1_168 ({gpcOutL0_193[0], gpcOutL0_192[1], gpcOutL0_191[2], gpcOutL0_89[0], gpcOutL0_88[1], gpcOutL0_87[2]}, gpcOutL1_168);
gpc006 gpcL1_169 ({gpcOutL0_194[0], gpcOutL0_193[1], gpcOutL0_192[2], gpcOutL0_90[0], gpcOutL0_89[1], gpcOutL0_88[2]}, gpcOutL1_169);
gpc006 gpcL1_170 ({gpcOutL0_195[0], gpcOutL0_194[1], gpcOutL0_193[2], gpcOutL0_91[0], gpcOutL0_90[1], gpcOutL0_89[2]}, gpcOutL1_170);
gpc006 gpcL1_171 ({gpcOutL0_195[2], gpcOutL0_93[0], gpcOutL0_92[1], gpcOutL0_91[2], pp319[3], pp303[5]}, gpcOutL1_171);
gpc006 gpcL1_172 ({gpcOutL0_142[0], gpcOutL0_141[1], gpcOutL0_140[2], gpcOutL0_38[0], gpcOutL0_37[1], gpcOutL0_36[2]}, gpcOutL1_172);
gpc006 gpcL1_173 ({gpcOutL0_144[0], gpcOutL0_143[1], gpcOutL0_142[2], gpcOutL0_40[0], gpcOutL0_39[1], gpcOutL0_38[2]}, gpcOutL1_173);
gpc006 gpcL1_174 ({gpcOutL0_145[0], gpcOutL0_144[1], gpcOutL0_143[2], gpcOutL0_41[0], gpcOutL0_40[1], gpcOutL0_39[2]}, gpcOutL1_174);
gpc006 gpcL1_175 ({gpcOutL0_232[2], gpcOutL0_146[0], gpcOutL0_145[1], gpcOutL0_144[2], gpcOutL0_42[0], gpcOutL0_41[1]}, gpcOutL1_175);
gpc006 gpcL1_176 ({gpcOutL0_233[2], gpcOutL0_147[0], gpcOutL0_146[1], gpcOutL0_145[2], gpcOutL0_43[0], gpcOutL0_42[1]}, gpcOutL1_176);
gpc006 gpcL1_177 ({gpcOutL0_235[1], gpcOutL0_234[2], gpcOutL0_148[0], gpcOutL0_147[1], gpcOutL0_146[2], gpcOutL0_44[0]}, gpcOutL1_177);
gpc006 gpcL1_178 ({gpcOutL0_236[1], gpcOutL0_235[2], gpcOutL0_149[0], gpcOutL0_148[1], gpcOutL0_147[2], gpcOutL0_45[0]}, gpcOutL1_178);
gpc006 gpcL1_179 ({gpcOutL0_238[0], gpcOutL0_237[1], gpcOutL0_236[2], gpcOutL0_150[0], gpcOutL0_149[1], gpcOutL0_148[2]}, gpcOutL1_179);
gpc006 gpcL1_180 ({gpcOutL0_238[1], gpcOutL0_237[2], gpcOutL0_151[0], gpcOutL0_150[1], gpcOutL0_149[2], gpcOutL0_47[0]}, gpcOutL1_180);
gpc006 gpcL1_181 ({gpcOutL0_240[0], gpcOutL0_239[1], gpcOutL0_238[2], gpcOutL0_152[0], gpcOutL0_151[1], gpcOutL0_150[2]}, gpcOutL1_181);
gpc006 gpcL1_182 ({gpcOutL0_241[0], gpcOutL0_240[1], gpcOutL0_239[2], gpcOutL0_153[0], gpcOutL0_152[1], gpcOutL0_151[2]}, gpcOutL1_182);
gpc006 gpcL1_183 ({gpcOutL0_312[2], gpcOutL0_242[0], gpcOutL0_241[1], gpcOutL0_240[2], gpcOutL0_154[0], gpcOutL0_153[1]}, gpcOutL1_183);
gpc006 gpcL1_184 ({gpcOutL0_313[2], gpcOutL0_243[0], gpcOutL0_242[1], gpcOutL0_241[2], gpcOutL0_155[0], gpcOutL0_154[1]}, gpcOutL1_184);
gpc006 gpcL1_185 ({gpcOutL0_315[1], gpcOutL0_314[2], gpcOutL0_244[0], gpcOutL0_243[1], gpcOutL0_242[2], gpcOutL0_156[0]}, gpcOutL1_185);
gpc006 gpcL1_186 ({gpcOutL0_316[1], gpcOutL0_315[2], gpcOutL0_245[0], gpcOutL0_244[1], gpcOutL0_243[2], gpcOutL0_157[0]}, gpcOutL1_186);
gpc006 gpcL1_187 ({gpcOutL0_318[0], gpcOutL0_317[1], gpcOutL0_316[2], gpcOutL0_246[0], gpcOutL0_245[1], gpcOutL0_244[2]}, gpcOutL1_187);
gpc006 gpcL1_188 ({gpcOutL0_318[1], gpcOutL0_317[2], gpcOutL0_247[0], gpcOutL0_246[1], gpcOutL0_245[2], gpcOutL0_159[0]}, gpcOutL1_188);
gpc006 gpcL1_189 ({gpcOutL0_320[0], gpcOutL0_319[1], gpcOutL0_318[2], gpcOutL0_248[0], gpcOutL0_247[1], gpcOutL0_246[2]}, gpcOutL1_189);
gpc006 gpcL1_190 ({gpcOutL0_320[1], gpcOutL0_319[2], gpcOutL0_249[0], gpcOutL0_248[1], gpcOutL0_247[2], gpcOutL0_161[0]}, gpcOutL1_190);
gpc006 gpcL1_191 ({gpcOutL0_322[0], gpcOutL0_321[1], gpcOutL0_320[2], gpcOutL0_250[0], gpcOutL0_249[1], gpcOutL0_248[2]}, gpcOutL1_191);
gpc006 gpcL1_192 ({gpcOutL0_323[0], gpcOutL0_322[1], gpcOutL0_321[2], gpcOutL0_251[0], gpcOutL0_250[1], gpcOutL0_249[2]}, gpcOutL1_192);
gpc006 gpcL1_193 ({gpcOutL0_322[2], gpcOutL0_252[0], gpcOutL0_251[1], gpcOutL0_250[2], gpcOutL0_164[0], gpcOutL0_163[1]}, gpcOutL1_193);
gpc006 gpcL1_194 ({gpcOutL0_323[2], gpcOutL0_253[0], gpcOutL0_252[1], gpcOutL0_251[2], gpcOutL0_165[0], gpcOutL0_164[1]}, gpcOutL1_194);
gpc006 gpcL1_195 ({gpcOutL0_254[0], gpcOutL0_253[1], gpcOutL0_252[2], gpcOutL0_166[0], gpcOutL0_165[1], gpcOutL0_164[2]}, gpcOutL1_195);
gpc006 gpcL1_196 ({gpcOutL0_255[0], gpcOutL0_254[1], gpcOutL0_253[2], gpcOutL0_167[0], gpcOutL0_166[1], gpcOutL0_165[2]}, gpcOutL1_196);
gpc006 gpcL1_197 ({gpcOutL0_256[0], gpcOutL0_255[1], gpcOutL0_254[2], gpcOutL0_168[0], gpcOutL0_167[1], gpcOutL0_166[2]}, gpcOutL1_197);
gpc006 gpcL1_198 ({gpcOutL0_257[0], gpcOutL0_256[1], gpcOutL0_255[2], gpcOutL0_169[0], gpcOutL0_168[1], gpcOutL0_167[2]}, gpcOutL1_198);
gpc006 gpcL1_199 ({gpcOutL0_258[0], gpcOutL0_257[1], gpcOutL0_256[2], gpcOutL0_170[0], gpcOutL0_169[1], gpcOutL0_168[2]}, gpcOutL1_199);
gpc006 gpcL1_200 ({gpcOutL0_259[0], gpcOutL0_258[1], gpcOutL0_257[2], gpcOutL0_171[0], gpcOutL0_170[1], gpcOutL0_169[2]}, gpcOutL1_200);
gpc006 gpcL1_201 ({gpcOutL0_258[2], gpcOutL0_172[0], gpcOutL0_171[1], gpcOutL0_170[2], gpcOutL0_68[0], gpcOutL0_67[1]}, gpcOutL1_201);
gpc006 gpcL1_202 ({gpcOutL0_259[2], gpcOutL0_173[0], gpcOutL0_172[1], gpcOutL0_171[2], gpcOutL0_69[0], gpcOutL0_68[1]}, gpcOutL1_202);
gpc006 gpcL1_203 ({gpcOutL0_174[0], gpcOutL0_173[1], gpcOutL0_172[2], gpcOutL0_70[0], gpcOutL0_69[1], gpcOutL0_68[2]}, gpcOutL1_203);
gpc006 gpcL1_204 ({gpcOutL0_175[0], gpcOutL0_174[1], gpcOutL0_173[2], gpcOutL0_71[0], gpcOutL0_70[1], gpcOutL0_69[2]}, gpcOutL1_204);
gpc006 gpcL1_205 ({gpcOutL0_176[0], gpcOutL0_175[1], gpcOutL0_174[2], gpcOutL0_72[0], gpcOutL0_71[1], gpcOutL0_70[2]}, gpcOutL1_205);
gpc006 gpcL1_206 ({gpcOutL0_177[0], gpcOutL0_176[1], gpcOutL0_175[2], gpcOutL0_73[0], gpcOutL0_72[1], gpcOutL0_71[2]}, gpcOutL1_206);
gpc006 gpcL1_207 ({gpcOutL0_178[0], gpcOutL0_177[1], gpcOutL0_176[2], gpcOutL0_74[0], gpcOutL0_73[1], gpcOutL0_72[2]}, gpcOutL1_207);
gpc006 gpcL1_208 ({gpcOutL0_179[0], gpcOutL0_178[1], gpcOutL0_177[2], gpcOutL0_75[0], gpcOutL0_74[1], gpcOutL0_73[2]}, gpcOutL1_208);
gpc006 gpcL1_209 ({gpcOutL0_179[2], gpcOutL0_77[0], gpcOutL0_76[1], gpcOutL0_75[2], pp191[3], pp175[5]}, gpcOutL1_209);
gpc006 gpcL1_210 ({gpcOutL0_158[0], gpcOutL0_157[1], gpcOutL0_156[2], gpcOutL0_54[0], gpcOutL0_53[1], gpcOutL0_52[2]}, gpcOutL1_210);
gpc006 gpcL1_211 ({gpcOutL0_158[1], gpcOutL0_157[2], gpcOutL0_55[0], gpcOutL0_54[1], gpcOutL0_53[2], pp15[3]}, gpcOutL1_211);
gpc006 gpcL1_212 ({gpcOutL0_160[0], gpcOutL0_159[1], gpcOutL0_158[2], gpcOutL0_56[0], gpcOutL0_55[1], gpcOutL0_54[2]}, gpcOutL1_212);
gpc006 gpcL1_213 ({gpcOutL0_162[0], gpcOutL0_161[1], gpcOutL0_160[2], gpcOutL0_58[0], gpcOutL0_57[1], gpcOutL0_56[2]}, gpcOutL1_213);
gpc006 gpcL1_214 ({gpcOutL0_163[0], gpcOutL0_162[1], gpcOutL0_161[2], gpcOutL0_59[0], gpcOutL0_58[1], gpcOutL0_57[2]}, gpcOutL1_214);
gpc006 gpcL1_215 ({gpcOutL0_163[2], gpcOutL0_61[0], gpcOutL0_60[1], gpcOutL0_59[2], pp63[3], pp47[5]}, gpcOutL1_215);
gpc015 gpcL1_216 ({gpcOutL0_496[0], gpcOutL0_512[2], gpcOutL0_466[0], gpcOutL0_4[0], gpcOutL0_3[1], gpcOutL0_2[2]}, gpcOutL1_216);
gpc015 gpcL1_217 ({gpcOutL0_124[1], gpcOutL0_123[1], gpcOutL0_122[2], gpcOutL0_20[0], gpcOutL0_19[1], gpcOutL0_18[2]}, gpcOutL1_217);
gpc015 gpcL1_218 ({gpcOutL0_140[1], gpcOutL0_139[1], gpcOutL0_138[2], gpcOutL0_36[0], gpcOutL0_35[1], gpcOutL0_34[2]}, gpcOutL1_218);
gpc015 gpcL1_219 ({gpcOutL0_156[1], gpcOutL0_155[1], gpcOutL0_154[2], gpcOutL0_52[0], gpcOutL0_51[1], gpcOutL0_50[2]}, gpcOutL1_219);
gpc005 gpcL1_220 ({gpcOutL0_467[0], gpcOutL0_449[1], gpcOutL0_7[0], gpcOutL0_6[1], gpcOutL0_5[2]}, gpcOutL1_220);
gpc005 gpcL1_221 ({gpcOutL0_126[1], gpcOutL0_125[2], gpcOutL0_23[0], gpcOutL0_22[1], gpcOutL0_21[2]}, gpcOutL1_221);
gpc005 gpcL1_222 ({gpcOutL0_142[1], gpcOutL0_141[2], gpcOutL0_39[0], gpcOutL0_38[1], gpcOutL0_37[2]}, gpcOutL1_222);
gpc005 gpcL1_223 ({gpcOutL0_160[1], gpcOutL0_159[2], gpcOutL0_57[0], gpcOutL0_56[1], gpcOutL0_55[2]}, gpcOutL1_223);
gpc005 gpcL1_224 ({gpcOutL0_162[2], gpcOutL0_60[0], gpcOutL0_59[1], gpcOutL0_58[2], pp47[4]}, gpcOutL1_224);
gpc005 gpcL1_225 ({gpcOutL0_178[2], gpcOutL0_76[0], gpcOutL0_75[1], gpcOutL0_74[2], pp175[4]}, gpcOutL1_225);
gpc005 gpcL1_226 ({gpcOutL0_194[2], gpcOutL0_92[0], gpcOutL0_91[1], gpcOutL0_90[2], pp303[4]}, gpcOutL1_226);
gpc005 gpcL1_227 ({gpcOutL0_492[1], gpcOutL0_108[0], gpcOutL0_107[1], gpcOutL0_106[2], pp431[4]}, gpcOutL1_227);
gpc014 gpcL1_228 ({gpcOutL0_512[0], gpcOutL0_465[2], gpcOutL0_1[0], gpcOutL0_0[1], pp1[5]}, gpcOutL1_228);
gpc014 gpcL1_229 ({gpcOutL0_120[2], gpcOutL0_17[0], gpcOutL0_16[1], gpcOutL0_15[2], pp5[5]}, gpcOutL1_229);
gpc014 gpcL1_230 ({gpcOutL0_136[2], gpcOutL0_33[0], gpcOutL0_32[1], gpcOutL0_31[2], pp9[5]}, gpcOutL1_230);
gpc014 gpcL1_231 ({gpcOutL0_152[2], gpcOutL0_49[0], gpcOutL0_48[1], gpcOutL0_47[2], pp13[5]}, gpcOutL1_231);
gpc014 gpcL1_232 ({gpcOutL0_63[0], gpcOutL0_62[0], gpcOutL0_61[1], gpcOutL0_60[2], pp63[4]}, gpcOutL1_232);
gpc014 gpcL1_233 ({gpcOutL0_79[0], gpcOutL0_78[0], gpcOutL0_77[1], gpcOutL0_76[2], pp191[4]}, gpcOutL1_233);
gpc014 gpcL1_234 ({gpcOutL0_95[0], gpcOutL0_94[0], gpcOutL0_93[1], gpcOutL0_92[2], pp319[4]}, gpcOutL1_234);
gpc014 gpcL1_235 ({gpcOutL0_111[0], gpcOutL0_110[0], gpcOutL0_109[1], gpcOutL0_108[2], pp447[4]}, gpcOutL1_235);
gpc023 gpcL1_236 ({gpcOutL0_512[1], gpcOutL0_3[0], gpcOutL0_2[0], gpcOutL0_1[1], gpcOutL0_0[2]}, gpcOutL1_236);
gpc023 gpcL1_237 ({gpcOutL0_14[1], gpcOutL0_13[2], gpcOutL0_14[0], gpcOutL0_13[1], gpcOutL0_12[2]}, gpcOutL1_237);
gpc023 gpcL1_238 ({gpcOutL0_121[2], gpcOutL0_19[0], gpcOutL0_18[0], gpcOutL0_17[1], gpcOutL0_16[2]}, gpcOutL1_238);
gpc023 gpcL1_239 ({gpcOutL0_30[1], gpcOutL0_29[2], gpcOutL0_30[0], gpcOutL0_29[1], gpcOutL0_28[2]}, gpcOutL1_239);
gpc023 gpcL1_240 ({gpcOutL0_137[2], gpcOutL0_35[0], gpcOutL0_34[0], gpcOutL0_33[1], gpcOutL0_32[2]}, gpcOutL1_240);
gpc023 gpcL1_241 ({gpcOutL0_46[1], gpcOutL0_45[2], gpcOutL0_46[0], gpcOutL0_45[1], gpcOutL0_44[2]}, gpcOutL1_241);
gpc023 gpcL1_242 ({gpcOutL0_153[2], gpcOutL0_51[0], gpcOutL0_50[0], gpcOutL0_49[1], gpcOutL0_48[2]}, gpcOutL1_242);
gpc023 gpcL1_243 ({gpcOutL0_64[0], gpcOutL0_63[1], gpcOutL0_62[1], gpcOutL0_61[2], pp63[5]}, gpcOutL1_243);
gpc023 gpcL1_244 ({gpcOutL0_66[0], gpcOutL0_65[1], gpcOutL0_65[0], gpcOutL0_64[1], gpcOutL0_63[2]}, gpcOutL1_244);
gpc023 gpcL1_245 ({gpcOutL0_66[2], pp111[4], gpcOutL0_67[0], gpcOutL0_66[1], gpcOutL0_65[2]}, gpcOutL1_245);
gpc023 gpcL1_246 ({gpcOutL0_80[0], gpcOutL0_79[1], gpcOutL0_78[1], gpcOutL0_77[2], pp191[5]}, gpcOutL1_246);
gpc023 gpcL1_247 ({gpcOutL0_82[0], gpcOutL0_81[1], gpcOutL0_81[0], gpcOutL0_80[1], gpcOutL0_79[2]}, gpcOutL1_247);
gpc023 gpcL1_248 ({gpcOutL0_82[2], pp239[4], gpcOutL0_83[0], gpcOutL0_82[1], gpcOutL0_81[2]}, gpcOutL1_248);
gpc023 gpcL1_249 ({gpcOutL0_96[0], gpcOutL0_95[1], gpcOutL0_94[1], gpcOutL0_93[2], pp319[5]}, gpcOutL1_249);
gpc023 gpcL1_250 ({gpcOutL0_98[0], gpcOutL0_97[1], gpcOutL0_97[0], gpcOutL0_96[1], gpcOutL0_95[2]}, gpcOutL1_250);
gpc023 gpcL1_251 ({gpcOutL0_98[2], pp367[4], gpcOutL0_99[0], gpcOutL0_98[1], gpcOutL0_97[2]}, gpcOutL1_251);
gpc023 gpcL1_252 ({gpcOutL0_463[0], gpcOutL0_111[1], gpcOutL0_110[1], gpcOutL0_109[2], pp447[5]}, gpcOutL1_252);
gpc023 gpcL1_253 ({gpcOutL0_511[0], gpcOutL0_493[1], gpcOutL0_493[0], gpcOutL0_463[1], gpcOutL0_111[2]}, gpcOutL1_253);
gpc023 gpcL1_254 ({gpcOutL0_494[1], pp495[4], gpcOutL0_511[1], gpcOutL0_494[0], gpcOutL0_493[2]}, gpcOutL1_254);
gpc003 gpcL1_255 ({gpcOutL0_466[1], gpcOutL0_5[0], gpcOutL0_4[1]}, gpcOutL1_255);
gpc003 gpcL1_256 ({gpcOutL0_16[0], gpcOutL0_15[1], gpcOutL0_14[2]}, gpcOutL1_256);
gpc003 gpcL1_257 ({gpcOutL0_123[2], gpcOutL0_21[0], gpcOutL0_20[1]}, gpcOutL1_257);
gpc003 gpcL1_258 ({gpcOutL0_32[0], gpcOutL0_31[1], gpcOutL0_30[2]}, gpcOutL1_258);
gpc003 gpcL1_259 ({gpcOutL0_139[2], gpcOutL0_37[0], gpcOutL0_36[1]}, gpcOutL1_259);
gpc003 gpcL1_260 ({gpcOutL0_48[0], gpcOutL0_47[1], gpcOutL0_46[2]}, gpcOutL1_260);
gpc003 gpcL1_261 ({gpcOutL0_155[2], gpcOutL0_53[0], gpcOutL0_52[1]}, gpcOutL1_261);
gpc003 gpcL1_262 ({gpcOutL0_67[2], pp127[3], pp111[5]}, gpcOutL1_262);
gpc003 gpcL1_263 ({gpcOutL0_83[2], pp255[3], pp239[5]}, gpcOutL1_263);
gpc003 gpcL1_264 ({gpcOutL0_99[2], pp383[3], pp367[5]}, gpcOutL1_264);
gpc003 gpcL1_265 ({gpcOutL0_494[2], pp511[3], pp495[5]}, gpcOutL1_265);
gpc022 gpcL1_266 ({gpcOutL0_12[1], gpcOutL0_11[2], gpcOutL0_11[1], gpcOutL0_10[2]}, gpcOutL1_266);
gpc022 gpcL1_267 ({gpcOutL0_28[1], gpcOutL0_27[2], gpcOutL0_27[1], gpcOutL0_26[2]}, gpcOutL1_267);
gpc022 gpcL1_268 ({gpcOutL0_44[1], gpcOutL0_43[2], gpcOutL0_43[1], gpcOutL0_42[2]}, gpcOutL1_268);
gpc222 gpcL1_269 ({gpcOutL0_495[1], gpcOutL0_464[2], gpcOutL0_495[0], gpcOutL0_464[1], gpcOutL0_519[2], gpcOutL0_464[0]}, gpcOutL1_269);

// level 2
wire [2:0]  gpcOutL2_0;
wire [2:0]  gpcOutL2_1;
wire [2:0]  gpcOutL2_2;
wire [2:0]  gpcOutL2_3;
wire [2:0]  gpcOutL2_4;
wire [2:0]  gpcOutL2_5;
wire [2:0]  gpcOutL2_6;
wire [2:0]  gpcOutL2_7;
wire [2:0]  gpcOutL2_8;
wire [2:0]  gpcOutL2_9;
wire [2:0]  gpcOutL2_10;
wire [2:0]  gpcOutL2_11;
wire [2:0]  gpcOutL2_12;
wire [2:0]  gpcOutL2_13;
wire [2:0]  gpcOutL2_14;
wire [2:0]  gpcOutL2_15;
wire [2:0]  gpcOutL2_16;
wire [2:0]  gpcOutL2_17;
wire [2:0]  gpcOutL2_18;
wire [2:0]  gpcOutL2_19;
wire [2:0]  gpcOutL2_20;
wire [2:0]  gpcOutL2_21;
wire [2:0]  gpcOutL2_22;
wire [2:0]  gpcOutL2_23;
wire [2:0]  gpcOutL2_24;
wire [2:0]  gpcOutL2_25;
wire [2:0]  gpcOutL2_26;
wire [2:0]  gpcOutL2_27;
wire [2:0]  gpcOutL2_28;
wire [2:0]  gpcOutL2_29;
wire [2:0]  gpcOutL2_30;
wire [2:0]  gpcOutL2_31;
wire [2:0]  gpcOutL2_32;
wire [2:0]  gpcOutL2_33;
wire [2:0]  gpcOutL2_34;
wire [2:0]  gpcOutL2_35;
wire [2:0]  gpcOutL2_36;
wire [2:0]  gpcOutL2_37;
wire [2:0]  gpcOutL2_38;
wire [2:0]  gpcOutL2_39;
wire [2:0]  gpcOutL2_40;
wire [2:0]  gpcOutL2_41;
wire [2:0]  gpcOutL2_42;
wire [2:0]  gpcOutL2_43;
wire [2:0]  gpcOutL2_44;
wire [2:0]  gpcOutL2_45;
wire [2:0]  gpcOutL2_46;
wire [2:0]  gpcOutL2_47;
wire [2:0]  gpcOutL2_48;
wire [2:0]  gpcOutL2_49;
wire [2:0]  gpcOutL2_50;
wire [2:0]  gpcOutL2_51;
wire [2:0]  gpcOutL2_52;
wire [2:0]  gpcOutL2_53;
wire [2:0]  gpcOutL2_54;
wire [2:0]  gpcOutL2_55;
wire [2:0]  gpcOutL2_56;
wire [2:0]  gpcOutL2_57;
wire [2:0]  gpcOutL2_58;
wire [2:0]  gpcOutL2_59;
wire [2:0]  gpcOutL2_60;
wire [2:0]  gpcOutL2_61;
wire [2:0]  gpcOutL2_62;
wire [2:0]  gpcOutL2_63;
wire [2:0]  gpcOutL2_64;
wire [2:0]  gpcOutL2_65;
wire [2:0]  gpcOutL2_66;
wire [2:0]  gpcOutL2_67;
wire [2:0]  gpcOutL2_68;
wire [2:0]  gpcOutL2_69;
wire [2:0]  gpcOutL2_70;
wire [2:0]  gpcOutL2_71;
wire [2:0]  gpcOutL2_72;
wire [2:0]  gpcOutL2_73;
wire [2:0]  gpcOutL2_74;
wire [2:0]  gpcOutL2_75;
wire [2:0]  gpcOutL2_76;
wire [2:0]  gpcOutL2_77;
wire [2:0]  gpcOutL2_78;
wire [2:0]  gpcOutL2_79;
wire [2:0]  gpcOutL2_80;
wire [2:0]  gpcOutL2_81;
wire [2:0]  gpcOutL2_82;
wire [2:0]  gpcOutL2_83;
wire [2:0]  gpcOutL2_84;
wire [2:0]  gpcOutL2_85;
wire [2:0]  gpcOutL2_86;
wire [2:0]  gpcOutL2_87;
wire [2:0]  gpcOutL2_88;
wire [2:0]  gpcOutL2_89;
wire [2:0]  gpcOutL2_90;
wire [2:0]  gpcOutL2_91;
wire [2:0]  gpcOutL2_92;
wire [2:0]  gpcOutL2_93;
wire [2:0]  gpcOutL2_94;
wire [2:0]  gpcOutL2_95;
wire [2:0]  gpcOutL2_96;
wire [2:0]  gpcOutL2_97;
wire [2:0]  gpcOutL2_98;
wire [2:0]  gpcOutL2_99;
wire [2:0]  gpcOutL2_100;
wire [2:0]  gpcOutL2_101;
wire [2:0]  gpcOutL2_102;
wire [2:0]  gpcOutL2_103;
wire [2:0]  gpcOutL2_104;
wire [2:0]  gpcOutL2_105;
wire [2:0]  gpcOutL2_106;
wire [2:0]  gpcOutL2_107;
wire [2:0]  gpcOutL2_108;
wire [2:0]  gpcOutL2_109;
wire [2:0]  gpcOutL2_110;
wire [2:0]  gpcOutL2_111;
wire [2:0]  gpcOutL2_112;
wire [2:0]  gpcOutL2_113;
wire [2:0]  gpcOutL2_114;
wire [2:0]  gpcOutL2_115;
wire [2:0]  gpcOutL2_116;
wire [2:0]  gpcOutL2_117;
wire [2:0]  gpcOutL2_118;
wire [2:0]  gpcOutL2_119;
wire [2:0]  gpcOutL2_120;
wire [2:0]  gpcOutL2_121;
wire [2:0]  gpcOutL2_122;
wire [2:0]  gpcOutL2_123;
wire [2:0]  gpcOutL2_124;
wire [2:0]  gpcOutL2_125;
wire [3:0]  gpcOutL2_126;
wire [3:0]  gpcOutL2_127;
wire [1:0]  gpcOutL2_128;
wire [1:0]  gpcOutL2_129;
wire [1:0]  gpcOutL2_130;
wire [1:0]  gpcOutL2_131;
wire [1:0]  gpcOutL2_132;
wire [1:0]  gpcOutL2_133;
wire [1:0]  gpcOutL2_134;
wire [1:0]  gpcOutL2_135;
wire [1:0]  gpcOutL2_136;
wire [1:0]  gpcOutL2_137;
wire [1:0]  gpcOutL2_138;
wire [2:0]  gpcOutL2_139;
wire [3:0]  gpcOutL2_140;

gpc006 gpcL2_0 ({gpcOutL1_238[1], gpcOutL1_229[2], gpcOutL1_12[0], gpcOutL1_11[1], gpcOutL1_10[2], gpcOutL0_18[1]}, gpcOutL2_0);
gpc006 gpcL2_1 ({gpcOutL1_257[0], gpcOutL1_217[1], gpcOutL1_14[0], gpcOutL1_13[1], gpcOutL1_12[2], gpcOutL0_19[2]}, gpcOutL2_1);
gpc006 gpcL2_2 ({gpcOutL1_257[1], gpcOutL1_217[2], gpcOutL1_102[0], gpcOutL1_15[0], gpcOutL1_14[1], gpcOutL1_13[2]}, gpcOutL2_2);
gpc006 gpcL2_3 ({gpcOutL1_221[1], gpcOutL1_103[0], gpcOutL1_102[2], gpcOutL1_17[0], gpcOutL1_16[1], gpcOutL1_15[2]}, gpcOutL2_3);
gpc006 gpcL2_4 ({gpcOutL1_221[2], gpcOutL1_104[0], gpcOutL1_103[1], gpcOutL1_18[0], gpcOutL1_17[1], gpcOutL1_16[2]}, gpcOutL2_4);
gpc006 gpcL2_5 ({gpcOutL1_105[0], gpcOutL1_104[1], gpcOutL1_103[2], gpcOutL1_19[0], gpcOutL1_18[1], gpcOutL1_17[2]}, gpcOutL2_5);
gpc006 gpcL2_6 ({gpcOutL1_106[0], gpcOutL1_105[1], gpcOutL1_104[2], gpcOutL1_20[0], gpcOutL1_19[1], gpcOutL1_18[2]}, gpcOutL2_6);
gpc006 gpcL2_7 ({gpcOutL1_267[0], gpcOutL1_107[0], gpcOutL1_106[1], gpcOutL1_105[2], gpcOutL1_21[0], gpcOutL1_20[1]}, gpcOutL2_7);
gpc006 gpcL2_8 ({gpcOutL1_267[1], gpcOutL1_108[0], gpcOutL1_107[1], gpcOutL1_106[2], gpcOutL1_22[0], gpcOutL1_21[1]}, gpcOutL2_8);
gpc006 gpcL2_9 ({gpcOutL1_267[2], gpcOutL1_239[0], gpcOutL1_109[0], gpcOutL1_108[1], gpcOutL1_107[2], gpcOutL1_23[0]}, gpcOutL2_9);
gpc006 gpcL2_10 ({gpcOutL1_239[1], gpcOutL1_110[0], gpcOutL1_109[1], gpcOutL1_108[2], gpcOutL1_24[0], gpcOutL1_23[1]}, gpcOutL2_10);
gpc006 gpcL2_11 ({gpcOutL1_258[0], gpcOutL1_239[2], gpcOutL1_111[0], gpcOutL1_110[1], gpcOutL1_109[2], gpcOutL1_25[0]}, gpcOutL2_11);
gpc006 gpcL2_12 ({gpcOutL1_258[1], gpcOutL1_230[0], gpcOutL1_112[0], gpcOutL1_111[1], gpcOutL1_110[2], gpcOutL1_26[0]}, gpcOutL2_12);
gpc006 gpcL2_13 ({gpcOutL1_240[0], gpcOutL1_230[1], gpcOutL1_113[0], gpcOutL1_112[1], gpcOutL1_111[2], gpcOutL1_27[0]}, gpcOutL2_13);
gpc006 gpcL2_14 ({gpcOutL1_240[1], gpcOutL1_230[2], gpcOutL1_114[0], gpcOutL1_113[1], gpcOutL1_112[2], gpcOutL1_28[0]}, gpcOutL2_14);
gpc006 gpcL2_15 ({gpcOutL1_240[2], gpcOutL1_218[0], gpcOutL1_115[0], gpcOutL1_114[1], gpcOutL1_113[2], gpcOutL1_29[0]}, gpcOutL2_15);
gpc006 gpcL2_16 ({gpcOutL1_259[0], gpcOutL1_218[1], gpcOutL1_116[0], gpcOutL1_115[1], gpcOutL1_114[2], gpcOutL1_30[0]}, gpcOutL2_16);
gpc006 gpcL2_17 ({gpcOutL1_259[1], gpcOutL1_218[2], gpcOutL1_172[0], gpcOutL1_117[0], gpcOutL1_116[1], gpcOutL1_115[2]}, gpcOutL2_17);
gpc006 gpcL2_18 ({gpcOutL1_222[0], gpcOutL1_172[1], gpcOutL1_118[0], gpcOutL1_117[1], gpcOutL1_116[2], gpcOutL1_32[0]}, gpcOutL2_18);
gpc006 gpcL2_19 ({gpcOutL1_222[1], gpcOutL1_173[0], gpcOutL1_172[2], gpcOutL1_119[0], gpcOutL1_118[1], gpcOutL1_117[2]}, gpcOutL2_19);
gpc006 gpcL2_20 ({gpcOutL1_222[2], gpcOutL1_174[0], gpcOutL1_173[1], gpcOutL1_120[0], gpcOutL1_119[1], gpcOutL1_118[2]}, gpcOutL2_20);
gpc006 gpcL2_21 ({gpcOutL1_175[0], gpcOutL1_174[1], gpcOutL1_173[2], gpcOutL1_121[0], gpcOutL1_120[1], gpcOutL1_119[2]}, gpcOutL2_21);
gpc006 gpcL2_22 ({gpcOutL1_176[0], gpcOutL1_175[1], gpcOutL1_174[2], gpcOutL1_122[0], gpcOutL1_121[1], gpcOutL1_120[2]}, gpcOutL2_22);
gpc006 gpcL2_23 ({gpcOutL1_268[0], gpcOutL1_177[0], gpcOutL1_176[1], gpcOutL1_175[2], gpcOutL1_123[0], gpcOutL1_122[1]}, gpcOutL2_23);
gpc006 gpcL2_24 ({gpcOutL1_268[1], gpcOutL1_178[0], gpcOutL1_177[1], gpcOutL1_176[2], gpcOutL1_124[0], gpcOutL1_123[1]}, gpcOutL2_24);
gpc006 gpcL2_25 ({gpcOutL1_268[2], gpcOutL1_241[0], gpcOutL1_179[0], gpcOutL1_178[1], gpcOutL1_177[2], gpcOutL1_125[0]}, gpcOutL2_25);
gpc006 gpcL2_26 ({gpcOutL1_241[1], gpcOutL1_180[0], gpcOutL1_179[1], gpcOutL1_178[2], gpcOutL1_126[0], gpcOutL1_125[1]}, gpcOutL2_26);
gpc006 gpcL2_27 ({gpcOutL1_260[0], gpcOutL1_241[2], gpcOutL1_181[0], gpcOutL1_180[1], gpcOutL1_179[2], gpcOutL1_127[0]}, gpcOutL2_27);
gpc006 gpcL2_28 ({gpcOutL1_260[1], gpcOutL1_231[0], gpcOutL1_182[0], gpcOutL1_181[1], gpcOutL1_180[2], gpcOutL1_128[0]}, gpcOutL2_28);
gpc006 gpcL2_29 ({gpcOutL1_242[0], gpcOutL1_231[1], gpcOutL1_183[0], gpcOutL1_182[1], gpcOutL1_181[2], gpcOutL1_129[0]}, gpcOutL2_29);
gpc006 gpcL2_30 ({gpcOutL1_242[1], gpcOutL1_231[2], gpcOutL1_184[0], gpcOutL1_183[1], gpcOutL1_182[2], gpcOutL1_130[0]}, gpcOutL2_30);
gpc006 gpcL2_31 ({gpcOutL1_242[2], gpcOutL1_219[0], gpcOutL1_185[0], gpcOutL1_184[1], gpcOutL1_183[2], gpcOutL1_131[0]}, gpcOutL2_31);
gpc006 gpcL2_32 ({gpcOutL1_261[0], gpcOutL1_219[1], gpcOutL1_186[0], gpcOutL1_185[1], gpcOutL1_184[2], gpcOutL1_132[0]}, gpcOutL2_32);
gpc006 gpcL2_33 ({gpcOutL1_261[1], gpcOutL1_219[2], gpcOutL1_210[0], gpcOutL1_187[0], gpcOutL1_186[1], gpcOutL1_185[2]}, gpcOutL2_33);
gpc006 gpcL2_34 ({gpcOutL1_211[0], gpcOutL1_210[1], gpcOutL1_188[0], gpcOutL1_187[1], gpcOutL1_186[2], gpcOutL1_134[0]}, gpcOutL2_34);
gpc006 gpcL2_35 ({gpcOutL1_212[0], gpcOutL1_211[1], gpcOutL1_210[2], gpcOutL1_189[0], gpcOutL1_188[1], gpcOutL1_187[2]}, gpcOutL2_35);
gpc006 gpcL2_36 ({gpcOutL1_223[0], gpcOutL1_212[1], gpcOutL1_211[2], gpcOutL1_190[0], gpcOutL1_189[1], gpcOutL1_188[2]}, gpcOutL2_36);
gpc006 gpcL2_37 ({gpcOutL1_223[1], gpcOutL1_213[0], gpcOutL1_212[2], gpcOutL1_191[0], gpcOutL1_190[1], gpcOutL1_189[2]}, gpcOutL2_37);
gpc006 gpcL2_38 ({gpcOutL1_223[2], gpcOutL1_214[0], gpcOutL1_213[1], gpcOutL1_192[0], gpcOutL1_191[1], gpcOutL1_190[2]}, gpcOutL2_38);
gpc006 gpcL2_39 ({gpcOutL1_224[0], gpcOutL1_214[1], gpcOutL1_213[2], gpcOutL1_193[0], gpcOutL1_192[1], gpcOutL1_191[2]}, gpcOutL2_39);
gpc006 gpcL2_40 ({gpcOutL1_224[1], gpcOutL1_215[0], gpcOutL1_214[2], gpcOutL1_194[0], gpcOutL1_193[1], gpcOutL1_192[2]}, gpcOutL2_40);
gpc006 gpcL2_41 ({gpcOutL1_232[0], gpcOutL1_224[2], gpcOutL1_215[1], gpcOutL1_195[0], gpcOutL1_194[1], gpcOutL1_193[2]}, gpcOutL2_41);
gpc006 gpcL2_42 ({gpcOutL1_243[0], gpcOutL1_232[1], gpcOutL1_215[2], gpcOutL1_196[0], gpcOutL1_195[1], gpcOutL1_194[2]}, gpcOutL2_42);
gpc006 gpcL2_43 ({gpcOutL1_243[1], gpcOutL1_232[2], gpcOutL1_197[0], gpcOutL1_196[1], gpcOutL1_195[2], gpcOutL1_143[0]}, gpcOutL2_43);
gpc006 gpcL2_44 ({gpcOutL1_244[0], gpcOutL1_243[2], gpcOutL1_198[0], gpcOutL1_197[1], gpcOutL1_196[2], gpcOutL1_144[0]}, gpcOutL2_44);
gpc006 gpcL2_45 ({gpcOutL1_244[1], gpcOutL1_199[0], gpcOutL1_198[1], gpcOutL1_197[2], gpcOutL1_145[0], gpcOutL1_144[1]}, gpcOutL2_45);
gpc006 gpcL2_46 ({gpcOutL1_245[0], gpcOutL1_244[2], gpcOutL1_200[0], gpcOutL1_199[1], gpcOutL1_198[2], gpcOutL1_146[0]}, gpcOutL2_46);
gpc006 gpcL2_47 ({gpcOutL1_245[1], gpcOutL1_201[0], gpcOutL1_200[1], gpcOutL1_199[2], gpcOutL1_147[0], gpcOutL1_146[1]}, gpcOutL2_47);
gpc006 gpcL2_48 ({gpcOutL1_262[0], gpcOutL1_245[2], gpcOutL1_202[0], gpcOutL1_201[1], gpcOutL1_200[2], gpcOutL1_148[0]}, gpcOutL2_48);
gpc006 gpcL2_49 ({gpcOutL1_262[1], gpcOutL1_203[0], gpcOutL1_202[1], gpcOutL1_201[2], gpcOutL1_149[0], gpcOutL1_148[1]}, gpcOutL2_49);
gpc006 gpcL2_50 ({gpcOutL1_204[0], gpcOutL1_203[1], gpcOutL1_202[2], gpcOutL1_150[0], gpcOutL1_149[1], gpcOutL1_148[2]}, gpcOutL2_50);
gpc006 gpcL2_51 ({gpcOutL1_205[0], gpcOutL1_204[1], gpcOutL1_203[2], gpcOutL1_151[0], gpcOutL1_150[1], gpcOutL1_149[2]}, gpcOutL2_51);
gpc006 gpcL2_52 ({gpcOutL1_206[0], gpcOutL1_205[1], gpcOutL1_204[2], gpcOutL1_152[0], gpcOutL1_151[1], gpcOutL1_150[2]}, gpcOutL2_52);
gpc006 gpcL2_53 ({gpcOutL1_207[0], gpcOutL1_206[1], gpcOutL1_205[2], gpcOutL1_153[0], gpcOutL1_152[1], gpcOutL1_151[2]}, gpcOutL2_53);
gpc006 gpcL2_54 ({gpcOutL1_208[0], gpcOutL1_207[1], gpcOutL1_206[2], gpcOutL1_154[0], gpcOutL1_153[1], gpcOutL1_152[2]}, gpcOutL2_54);
gpc006 gpcL2_55 ({gpcOutL1_225[0], gpcOutL1_208[1], gpcOutL1_207[2], gpcOutL1_155[0], gpcOutL1_154[1], gpcOutL1_153[2]}, gpcOutL2_55);
gpc006 gpcL2_56 ({gpcOutL1_225[1], gpcOutL1_209[0], gpcOutL1_208[2], gpcOutL1_156[0], gpcOutL1_155[1], gpcOutL1_154[2]}, gpcOutL2_56);
gpc006 gpcL2_57 ({gpcOutL1_233[0], gpcOutL1_225[2], gpcOutL1_209[1], gpcOutL1_157[0], gpcOutL1_156[1], gpcOutL1_155[2]}, gpcOutL2_57);
gpc006 gpcL2_58 ({gpcOutL1_246[0], gpcOutL1_233[1], gpcOutL1_209[2], gpcOutL1_158[0], gpcOutL1_157[1], gpcOutL1_156[2]}, gpcOutL2_58);
gpc006 gpcL2_59 ({gpcOutL1_246[1], gpcOutL1_233[2], gpcOutL1_159[0], gpcOutL1_158[1], gpcOutL1_157[2], gpcOutL1_73[0]}, gpcOutL2_59);
gpc006 gpcL2_60 ({gpcOutL1_247[0], gpcOutL1_246[2], gpcOutL1_160[0], gpcOutL1_159[1], gpcOutL1_158[2], gpcOutL1_74[0]}, gpcOutL2_60);
gpc006 gpcL2_61 ({gpcOutL1_247[1], gpcOutL1_161[0], gpcOutL1_160[1], gpcOutL1_159[2], gpcOutL1_75[0], gpcOutL1_74[1]}, gpcOutL2_61);
gpc006 gpcL2_62 ({gpcOutL1_248[0], gpcOutL1_247[2], gpcOutL1_162[0], gpcOutL1_161[1], gpcOutL1_160[2], gpcOutL1_76[0]}, gpcOutL2_62);
gpc006 gpcL2_63 ({gpcOutL1_248[1], gpcOutL1_163[0], gpcOutL1_162[1], gpcOutL1_161[2], gpcOutL1_77[0], gpcOutL1_76[1]}, gpcOutL2_63);
gpc006 gpcL2_64 ({gpcOutL1_263[0], gpcOutL1_248[2], gpcOutL1_164[0], gpcOutL1_163[1], gpcOutL1_162[2], gpcOutL1_78[0]}, gpcOutL2_64);
gpc006 gpcL2_65 ({gpcOutL1_263[1], gpcOutL1_165[0], gpcOutL1_164[1], gpcOutL1_163[2], gpcOutL1_79[0], gpcOutL1_78[1]}, gpcOutL2_65);
gpc006 gpcL2_66 ({gpcOutL1_166[0], gpcOutL1_165[1], gpcOutL1_164[2], gpcOutL1_80[0], gpcOutL1_79[1], gpcOutL1_78[2]}, gpcOutL2_66);
gpc006 gpcL2_67 ({gpcOutL1_167[0], gpcOutL1_166[1], gpcOutL1_165[2], gpcOutL1_81[0], gpcOutL1_80[1], gpcOutL1_79[2]}, gpcOutL2_67);
gpc006 gpcL2_68 ({gpcOutL1_168[0], gpcOutL1_167[1], gpcOutL1_166[2], gpcOutL1_82[0], gpcOutL1_81[1], gpcOutL1_80[2]}, gpcOutL2_68);
gpc006 gpcL2_69 ({gpcOutL1_169[0], gpcOutL1_168[1], gpcOutL1_167[2], gpcOutL1_83[0], gpcOutL1_82[1], gpcOutL1_81[2]}, gpcOutL2_69);
gpc006 gpcL2_70 ({gpcOutL1_170[0], gpcOutL1_169[1], gpcOutL1_168[2], gpcOutL1_84[0], gpcOutL1_83[1], gpcOutL1_82[2]}, gpcOutL2_70);
gpc006 gpcL2_71 ({gpcOutL1_226[0], gpcOutL1_170[1], gpcOutL1_169[2], gpcOutL1_85[0], gpcOutL1_84[1], gpcOutL1_83[2]}, gpcOutL2_71);
gpc006 gpcL2_72 ({gpcOutL1_226[1], gpcOutL1_171[0], gpcOutL1_170[2], gpcOutL1_86[0], gpcOutL1_85[1], gpcOutL1_84[2]}, gpcOutL2_72);
gpc006 gpcL2_73 ({gpcOutL1_234[0], gpcOutL1_226[2], gpcOutL1_171[1], gpcOutL1_87[0], gpcOutL1_86[1], gpcOutL1_85[2]}, gpcOutL2_73);
gpc006 gpcL2_74 ({gpcOutL1_249[0], gpcOutL1_234[1], gpcOutL1_171[2], gpcOutL1_88[0], gpcOutL1_87[1], gpcOutL1_86[2]}, gpcOutL2_74);
gpc006 gpcL2_75 ({gpcOutL1_249[1], gpcOutL1_234[2], gpcOutL1_89[0], gpcOutL1_88[1], gpcOutL1_87[2], gpcOutL0_94[2]}, gpcOutL2_75);
gpc006 gpcL2_76 ({gpcOutL1_129[1], gpcOutL1_128[2], gpcOutL1_44[0], gpcOutL1_43[1], gpcOutL1_42[2], gpcOutL0_50[1]}, gpcOutL2_76);
gpc006 gpcL2_77 ({gpcOutL1_131[1], gpcOutL1_130[2], gpcOutL1_46[0], gpcOutL1_45[1], gpcOutL1_44[2], gpcOutL0_51[2]}, gpcOutL2_77);
gpc006 gpcL2_78 ({gpcOutL1_133[0], gpcOutL1_132[1], gpcOutL1_131[2], gpcOutL1_47[0], gpcOutL1_46[1], gpcOutL1_45[2]}, gpcOutL2_78);
gpc006 gpcL2_79 ({gpcOutL1_135[0], gpcOutL1_134[1], gpcOutL1_133[2], gpcOutL1_49[0], gpcOutL1_48[1], gpcOutL1_47[2]}, gpcOutL2_79);
gpc006 gpcL2_80 ({gpcOutL1_136[0], gpcOutL1_135[1], gpcOutL1_134[2], gpcOutL1_50[0], gpcOutL1_49[1], gpcOutL1_48[2]}, gpcOutL2_80);
gpc006 gpcL2_81 ({gpcOutL1_137[0], gpcOutL1_136[1], gpcOutL1_135[2], gpcOutL1_51[0], gpcOutL1_50[1], gpcOutL1_49[2]}, gpcOutL2_81);
gpc006 gpcL2_82 ({gpcOutL1_138[0], gpcOutL1_137[1], gpcOutL1_136[2], gpcOutL1_52[0], gpcOutL1_51[1], gpcOutL1_50[2]}, gpcOutL2_82);
gpc006 gpcL2_83 ({gpcOutL1_139[0], gpcOutL1_138[1], gpcOutL1_137[2], gpcOutL1_53[0], gpcOutL1_52[1], gpcOutL1_51[2]}, gpcOutL2_83);
gpc006 gpcL2_84 ({gpcOutL1_140[0], gpcOutL1_139[1], gpcOutL1_138[2], gpcOutL1_54[0], gpcOutL1_53[1], gpcOutL1_52[2]}, gpcOutL2_84);
gpc006 gpcL2_85 ({gpcOutL1_141[0], gpcOutL1_140[1], gpcOutL1_139[2], gpcOutL1_55[0], gpcOutL1_54[1], gpcOutL1_53[2]}, gpcOutL2_85);
gpc006 gpcL2_86 ({gpcOutL1_142[0], gpcOutL1_141[1], gpcOutL1_140[2], gpcOutL1_56[0], gpcOutL1_55[1], gpcOutL1_54[2]}, gpcOutL2_86);
gpc006 gpcL2_87 ({gpcOutL1_142[1], gpcOutL1_141[2], gpcOutL1_57[0], gpcOutL1_56[1], gpcOutL1_55[2], gpcOutL0_62[2]}, gpcOutL2_87);
gpc015 gpcL2_88 ({gpcOutL1_237[1], gpcOutL1_266[2], gpcOutL1_237[0], gpcOutL1_7[0], gpcOutL1_6[1], gpcOutL1_5[2]}, gpcOutL2_88);
gpc015 gpcL2_89 ({gpcOutL1_256[1], gpcOutL1_256[0], gpcOutL1_237[2], gpcOutL1_9[0], gpcOutL1_8[1], gpcOutL1_7[2]}, gpcOutL2_89);
gpc015 gpcL2_90 ({gpcOutL0_17[2], gpcOutL1_238[0], gpcOutL1_229[1], gpcOutL1_11[0], gpcOutL1_10[1], gpcOutL1_9[2]}, gpcOutL2_90);
gpc015 gpcL2_91 ({gpcOutL1_124[2], gpcOutL1_124[1], gpcOutL1_123[2], gpcOutL1_39[0], gpcOutL1_38[1], gpcOutL1_37[2]}, gpcOutL2_91);
gpc015 gpcL2_92 ({gpcOutL1_127[1], gpcOutL1_126[1], gpcOutL1_125[2], gpcOutL1_41[0], gpcOutL1_40[1], gpcOutL1_39[2]}, gpcOutL2_92);
gpc015 gpcL2_93 ({gpcOutL0_49[2], gpcOutL1_128[1], gpcOutL1_127[2], gpcOutL1_43[0], gpcOutL1_42[1], gpcOutL1_41[2]}, gpcOutL2_93);
gpc015 gpcL2_94 ({gpcOutL1_143[2], gpcOutL1_143[1], gpcOutL1_142[2], gpcOutL1_58[0], gpcOutL1_57[1], gpcOutL1_56[2]}, gpcOutL2_94);
gpc015 gpcL2_95 ({gpcOutL1_145[2], gpcOutL1_145[1], gpcOutL1_144[2], gpcOutL1_60[0], gpcOutL1_59[1], gpcOutL1_58[2]}, gpcOutL2_95);
gpc015 gpcL2_96 ({gpcOutL1_147[2], gpcOutL1_147[1], gpcOutL1_146[2], gpcOutL1_62[0], gpcOutL1_61[1], gpcOutL1_60[2]}, gpcOutL2_96);
gpc015 gpcL2_97 ({gpcOutL1_250[1], gpcOutL1_250[0], gpcOutL1_249[2], gpcOutL1_90[0], gpcOutL1_89[1], gpcOutL1_88[2]}, gpcOutL2_97);
gpc015 gpcL2_98 ({gpcOutL1_251[1], gpcOutL1_251[0], gpcOutL1_250[2], gpcOutL1_92[0], gpcOutL1_91[1], gpcOutL1_90[2]}, gpcOutL2_98);
gpc015 gpcL2_99 ({gpcOutL1_264[1], gpcOutL1_264[0], gpcOutL1_251[2], gpcOutL1_94[0], gpcOutL1_93[1], gpcOutL1_92[2]}, gpcOutL2_99);
gpc005 gpcL2_100 ({gpcOutL1_238[2], gpcOutL1_217[0], gpcOutL1_13[0], gpcOutL1_12[1], gpcOutL1_11[2]}, gpcOutL2_100);
gpc005 gpcL2_101 ({gpcOutL1_221[0], gpcOutL1_102[1], gpcOutL1_16[0], gpcOutL1_15[1], gpcOutL1_14[2]}, gpcOutL2_101);
gpc005 gpcL2_102 ({gpcOutL1_130[1], gpcOutL1_129[2], gpcOutL1_45[0], gpcOutL1_44[1], gpcOutL1_43[2]}, gpcOutL2_102);
gpc005 gpcL2_103 ({gpcOutL1_133[1], gpcOutL1_132[2], gpcOutL1_48[0], gpcOutL1_47[1], gpcOutL1_46[2]}, gpcOutL2_103);
gpc014 gpcL2_104 ({gpcOutL1_236[2], gpcOutL1_236[1], gpcOutL1_228[2], gpcOutL0_2[1], gpcOutL0_1[2]}, gpcOutL2_104);
gpc014 gpcL2_105 ({gpcOutL1_3[0], gpcOutL1_220[2], gpcOutL1_2[0], gpcOutL1_1[1], pp3[5]}, gpcOutL2_105);
gpc014 gpcL2_106 ({gpcOutL1_266[0], gpcOutL1_4[0], gpcOutL1_3[1], gpcOutL1_2[2], gpcOutL0_9[2]}, gpcOutL2_106);
gpc014 gpcL2_107 ({gpcOutL1_28[1], gpcOutL1_27[1], gpcOutL1_26[2], gpcOutL0_34[1], gpcOutL0_33[2]}, gpcOutL2_107);
gpc014 gpcL2_108 ({gpcOutL1_35[0], gpcOutL1_34[0], gpcOutL1_33[1], gpcOutL1_32[2], pp11[5]}, gpcOutL2_108);
gpc014 gpcL2_109 ({gpcOutL1_121[2], gpcOutL1_36[0], gpcOutL1_35[1], gpcOutL1_34[2], gpcOutL0_41[2]}, gpcOutL2_109);
gpc014 gpcL2_110 ({gpcOutL1_64[0], gpcOutL1_63[0], gpcOutL1_62[1], gpcOutL1_61[2], pp127[4]}, gpcOutL2_110);
gpc014 gpcL2_111 ({gpcOutL1_96[0], gpcOutL1_95[0], gpcOutL1_94[1], gpcOutL1_93[2], pp383[4]}, gpcOutL2_111);
gpc023 gpcL2_112 ({gpcOutL1_255[1], gpcOutL1_216[2], gpcOutL1_255[0], gpcOutL1_216[1], gpcOutL0_3[2]}, gpcOutL2_112);
gpc023 gpcL2_113 ({gpcOutL1_266[1], gpcOutL1_6[0], gpcOutL1_5[0], gpcOutL1_4[1], gpcOutL1_3[2]}, gpcOutL2_113);
gpc023 gpcL2_114 ({gpcOutL1_31[0], gpcOutL1_30[1], gpcOutL1_29[1], gpcOutL1_28[2], gpcOutL0_35[2]}, gpcOutL2_114);
gpc023 gpcL2_115 ({gpcOutL1_122[2], gpcOutL1_38[0], gpcOutL1_37[0], gpcOutL1_36[1], gpcOutL1_35[2]}, gpcOutL2_115);
gpc023 gpcL2_116 ({gpcOutL1_65[0], gpcOutL1_64[1], gpcOutL1_63[1], gpcOutL1_62[2], pp127[5]}, gpcOutL2_116);
gpc023 gpcL2_117 ({gpcOutL1_67[0], gpcOutL1_66[1], gpcOutL1_66[0], gpcOutL1_65[1], gpcOutL1_64[2]}, gpcOutL2_117);
gpc023 gpcL2_118 ({gpcOutL1_69[0], gpcOutL1_68[1], gpcOutL1_68[0], gpcOutL1_67[1], gpcOutL1_66[2]}, gpcOutL2_118);
gpc023 gpcL2_119 ({gpcOutL1_71[0], gpcOutL1_70[1], gpcOutL1_70[0], gpcOutL1_69[1], gpcOutL1_68[2]}, gpcOutL2_119);
gpc023 gpcL2_120 ({gpcOutL1_72[1], gpcOutL1_71[2], gpcOutL1_72[0], gpcOutL1_71[1], gpcOutL1_70[2]}, gpcOutL2_120);
gpc023 gpcL2_121 ({gpcOutL1_97[0], gpcOutL1_96[1], gpcOutL1_95[1], gpcOutL1_94[2], pp383[5]}, gpcOutL2_121);
gpc023 gpcL2_122 ({gpcOutL1_99[0], gpcOutL1_98[1], gpcOutL1_98[0], gpcOutL1_97[1], gpcOutL1_96[2]}, gpcOutL2_122);
gpc023 gpcL2_123 ({gpcOutL1_227[0], gpcOutL1_100[1], gpcOutL1_100[0], gpcOutL1_99[1], gpcOutL1_98[2]}, gpcOutL2_123);
gpc023 gpcL2_124 ({gpcOutL1_235[0], gpcOutL1_227[2], gpcOutL1_227[1], gpcOutL1_101[0], gpcOutL1_100[2]}, gpcOutL2_124);
gpc023 gpcL2_125 ({gpcOutL1_252[1], gpcOutL1_235[2], gpcOutL1_252[0], gpcOutL1_235[1], gpcOutL1_101[2]}, gpcOutL2_125);
gpc222 gpcL2_126 ({gpcOutL1_26[1], gpcOutL1_25[2], gpcOutL1_25[1], gpcOutL1_24[2], gpcOutL1_24[1], gpcOutL1_23[2]}, gpcOutL2_126);
gpc222 gpcL2_127 ({gpcOutL1_75[1], gpcOutL1_74[2], gpcOutL1_73[2], gpcOutL0_80[2], gpcOutL1_73[1], gpcOutL1_72[2]}, gpcOutL2_127);
gpc003 gpcL2_128 ({gpcOutL1_2[1], gpcOutL1_1[2], gpcOutL0_8[2]}, gpcOutL2_128);
gpc003 gpcL2_129 ({gpcOutL1_8[0], gpcOutL1_7[1], gpcOutL1_6[2]}, gpcOutL2_129);
gpc003 gpcL2_130 ({gpcOutL1_229[0], gpcOutL1_10[0], gpcOutL1_9[1]}, gpcOutL2_130);
gpc003 gpcL2_131 ({gpcOutL1_33[0], gpcOutL1_32[1], gpcOutL1_31[2]}, gpcOutL2_131);
gpc003 gpcL2_132 ({gpcOutL1_34[1], gpcOutL1_33[2], gpcOutL0_40[2]}, gpcOutL2_132);
gpc003 gpcL2_133 ({gpcOutL1_40[0], gpcOutL1_39[1], gpcOutL1_38[2]}, gpcOutL2_133);
gpc003 gpcL2_134 ({gpcOutL1_126[2], gpcOutL1_42[0], gpcOutL1_41[1]}, gpcOutL2_134);
gpc003 gpcL2_135 ({gpcOutL1_59[0], gpcOutL1_58[1], gpcOutL1_57[2]}, gpcOutL2_135);
gpc003 gpcL2_136 ({gpcOutL1_61[0], gpcOutL1_60[1], gpcOutL1_59[2]}, gpcOutL2_136);
gpc003 gpcL2_137 ({gpcOutL1_91[0], gpcOutL1_90[1], gpcOutL1_89[2]}, gpcOutL2_137);
gpc003 gpcL2_138 ({gpcOutL1_93[0], gpcOutL1_92[1], gpcOutL1_91[2]}, gpcOutL2_138);
gpc022 gpcL2_139 ({gpcOutL1_77[2], pp255[4], gpcOutL1_77[1], gpcOutL1_76[2]}, gpcOutL2_139);
gpc132 gpcL2_140 ({gpcOutL0_465[1], gpcOutL1_269[3], gpcOutL0_465[0], gpcOutL0_448[1], gpcOutL1_269[2], gpcOutL0_448[0]}, gpcOutL2_140);

// level 3
wire [2:0]  gpcOutL3_0;
wire [2:0]  gpcOutL3_1;
wire [2:0]  gpcOutL3_2;
wire [2:0]  gpcOutL3_3;
wire [2:0]  gpcOutL3_4;
wire [2:0]  gpcOutL3_5;
wire [2:0]  gpcOutL3_6;
wire [2:0]  gpcOutL3_7;
wire [2:0]  gpcOutL3_8;
wire [2:0]  gpcOutL3_9;
wire [2:0]  gpcOutL3_10;
wire [2:0]  gpcOutL3_11;
wire [2:0]  gpcOutL3_12;
wire [2:0]  gpcOutL3_13;
wire [2:0]  gpcOutL3_14;
wire [2:0]  gpcOutL3_15;
wire [2:0]  gpcOutL3_16;
wire [2:0]  gpcOutL3_17;
wire [2:0]  gpcOutL3_18;
wire [2:0]  gpcOutL3_19;
wire [2:0]  gpcOutL3_20;
wire [2:0]  gpcOutL3_21;
wire [2:0]  gpcOutL3_22;
wire [2:0]  gpcOutL3_23;
wire [2:0]  gpcOutL3_24;
wire [2:0]  gpcOutL3_25;
wire [2:0]  gpcOutL3_26;
wire [2:0]  gpcOutL3_27;
wire [2:0]  gpcOutL3_28;
wire [2:0]  gpcOutL3_29;
wire [2:0]  gpcOutL3_30;
wire [2:0]  gpcOutL3_31;
wire [2:0]  gpcOutL3_32;
wire [2:0]  gpcOutL3_33;
wire [2:0]  gpcOutL3_34;
wire [2:0]  gpcOutL3_35;
wire [2:0]  gpcOutL3_36;
wire [2:0]  gpcOutL3_37;
wire [2:0]  gpcOutL3_38;
wire [2:0]  gpcOutL3_39;
wire [2:0]  gpcOutL3_40;
wire [2:0]  gpcOutL3_41;
wire [2:0]  gpcOutL3_42;
wire [2:0]  gpcOutL3_43;
wire [2:0]  gpcOutL3_44;
wire [2:0]  gpcOutL3_45;
wire [2:0]  gpcOutL3_46;
wire [2:0]  gpcOutL3_47;
wire [2:0]  gpcOutL3_48;
wire [2:0]  gpcOutL3_49;
wire [2:0]  gpcOutL3_50;
wire [2:0]  gpcOutL3_51;
wire [2:0]  gpcOutL3_52;
wire [2:0]  gpcOutL3_53;
wire [1:0]  gpcOutL3_54;
wire [1:0]  gpcOutL3_55;
wire [1:0]  gpcOutL3_56;
wire [1:0]  gpcOutL3_57;
wire [1:0]  gpcOutL3_58;
wire [1:0]  gpcOutL3_59;
wire [1:0]  gpcOutL3_60;
wire [1:0]  gpcOutL3_61;
wire [1:0]  gpcOutL3_62;
wire [1:0]  gpcOutL3_63;
wire [1:0]  gpcOutL3_64;
wire [1:0]  gpcOutL3_65;
wire [2:0]  gpcOutL3_66;

gpc006 gpcL3_0 ({gpcOutL2_114[2], gpcOutL2_18[0], gpcOutL2_17[1], gpcOutL2_16[2], gpcOutL1_31[1], gpcOutL1_30[2]}, gpcOutL3_0);
gpc006 gpcL3_1 ({gpcOutL2_132[1], gpcOutL2_109[0], gpcOutL2_108[2], gpcOutL2_22[0], gpcOutL2_21[1], gpcOutL2_20[2]}, gpcOutL3_1);
gpc006 gpcL3_2 ({gpcOutL2_115[1], gpcOutL2_109[2], gpcOutL2_24[0], gpcOutL2_23[1], gpcOutL2_22[2], gpcOutL1_37[1]}, gpcOutL3_2);
gpc006 gpcL3_3 ({gpcOutL2_133[1], gpcOutL2_92[0], gpcOutL2_91[2], gpcOutL2_27[0], gpcOutL2_26[1], gpcOutL2_25[2]}, gpcOutL3_3);
gpc006 gpcL3_4 ({gpcOutL2_134[0], gpcOutL2_92[1], gpcOutL2_28[0], gpcOutL2_27[1], gpcOutL2_26[2], gpcOutL1_40[2]}, gpcOutL3_4);
gpc006 gpcL3_5 ({gpcOutL2_134[1], gpcOutL2_93[0], gpcOutL2_92[2], gpcOutL2_29[0], gpcOutL2_28[1], gpcOutL2_27[2]}, gpcOutL3_5);
gpc006 gpcL3_6 ({gpcOutL2_102[0], gpcOutL2_93[2], gpcOutL2_76[1], gpcOutL2_31[0], gpcOutL2_30[1], gpcOutL2_29[2]}, gpcOutL3_6);
gpc006 gpcL3_7 ({gpcOutL2_102[1], gpcOutL2_77[0], gpcOutL2_76[2], gpcOutL2_32[0], gpcOutL2_31[1], gpcOutL2_30[2]}, gpcOutL3_7);
gpc006 gpcL3_8 ({gpcOutL2_102[2], gpcOutL2_78[0], gpcOutL2_77[1], gpcOutL2_33[0], gpcOutL2_32[1], gpcOutL2_31[2]}, gpcOutL3_8);
gpc006 gpcL3_9 ({gpcOutL2_103[0], gpcOutL2_78[1], gpcOutL2_77[2], gpcOutL2_34[0], gpcOutL2_33[1], gpcOutL2_32[2]}, gpcOutL3_9);
gpc006 gpcL3_10 ({gpcOutL2_103[1], gpcOutL2_79[0], gpcOutL2_78[2], gpcOutL2_35[0], gpcOutL2_34[1], gpcOutL2_33[2]}, gpcOutL3_10);
gpc006 gpcL3_11 ({gpcOutL2_103[2], gpcOutL2_80[0], gpcOutL2_79[1], gpcOutL2_36[0], gpcOutL2_35[1], gpcOutL2_34[2]}, gpcOutL3_11);
gpc006 gpcL3_12 ({gpcOutL2_81[0], gpcOutL2_80[1], gpcOutL2_79[2], gpcOutL2_37[0], gpcOutL2_36[1], gpcOutL2_35[2]}, gpcOutL3_12);
gpc006 gpcL3_13 ({gpcOutL2_82[0], gpcOutL2_81[1], gpcOutL2_80[2], gpcOutL2_38[0], gpcOutL2_37[1], gpcOutL2_36[2]}, gpcOutL3_13);
gpc006 gpcL3_14 ({gpcOutL2_83[0], gpcOutL2_82[1], gpcOutL2_81[2], gpcOutL2_39[0], gpcOutL2_38[1], gpcOutL2_37[2]}, gpcOutL3_14);
gpc006 gpcL3_15 ({gpcOutL2_84[0], gpcOutL2_83[1], gpcOutL2_82[2], gpcOutL2_40[0], gpcOutL2_39[1], gpcOutL2_38[2]}, gpcOutL3_15);
gpc006 gpcL3_16 ({gpcOutL2_85[0], gpcOutL2_84[1], gpcOutL2_83[2], gpcOutL2_41[0], gpcOutL2_40[1], gpcOutL2_39[2]}, gpcOutL3_16);
gpc006 gpcL3_17 ({gpcOutL2_86[0], gpcOutL2_85[1], gpcOutL2_84[2], gpcOutL2_42[0], gpcOutL2_41[1], gpcOutL2_40[2]}, gpcOutL3_17);
gpc006 gpcL3_18 ({gpcOutL2_87[0], gpcOutL2_86[1], gpcOutL2_85[2], gpcOutL2_43[0], gpcOutL2_42[1], gpcOutL2_41[2]}, gpcOutL3_18);
gpc006 gpcL3_19 ({gpcOutL2_94[0], gpcOutL2_87[1], gpcOutL2_86[2], gpcOutL2_44[0], gpcOutL2_43[1], gpcOutL2_42[2]}, gpcOutL3_19);
gpc006 gpcL3_20 ({gpcOutL2_135[0], gpcOutL2_94[1], gpcOutL2_87[2], gpcOutL2_45[0], gpcOutL2_44[1], gpcOutL2_43[2]}, gpcOutL3_20);
gpc006 gpcL3_21 ({gpcOutL2_135[1], gpcOutL2_95[0], gpcOutL2_94[2], gpcOutL2_46[0], gpcOutL2_45[1], gpcOutL2_44[2]}, gpcOutL3_21);
gpc006 gpcL3_22 ({gpcOutL2_136[1], gpcOutL2_96[0], gpcOutL2_95[2], gpcOutL2_48[0], gpcOutL2_47[1], gpcOutL2_46[2]}, gpcOutL3_22);
gpc006 gpcL3_23 ({gpcOutL2_116[0], gpcOutL2_110[1], gpcOutL2_96[2], gpcOutL2_50[0], gpcOutL2_49[1], gpcOutL2_48[2]}, gpcOutL3_23);
gpc006 gpcL3_24 ({gpcOutL2_116[1], gpcOutL2_110[2], gpcOutL2_51[0], gpcOutL2_50[1], gpcOutL2_49[2], gpcOutL1_63[2]}, gpcOutL3_24);
gpc015 gpcL3_25 ({gpcOutL2_10[0], gpcOutL2_9[0], gpcOutL2_8[1], gpcOutL2_7[2], gpcOutL1_22[1], gpcOutL1_21[2]}, gpcOutL3_25);
gpc015 gpcL3_26 ({gpcOutL2_107[1], gpcOutL2_126[3], gpcOutL2_107[0], gpcOutL2_14[0], gpcOutL2_13[1], gpcOutL2_12[2]}, gpcOutL3_26);
gpc015 gpcL3_27 ({gpcOutL2_114[1], gpcOutL2_114[0], gpcOutL2_107[2], gpcOutL2_16[0], gpcOutL2_15[1], gpcOutL2_14[2]}, gpcOutL3_27);
gpc015 gpcL3_28 ({gpcOutL2_132[0], gpcOutL2_131[1], gpcOutL2_108[0], gpcOutL2_20[0], gpcOutL2_19[1], gpcOutL2_18[2]}, gpcOutL3_28);
gpc015 gpcL3_29 ({gpcOutL1_36[2], gpcOutL2_115[0], gpcOutL2_109[1], gpcOutL2_23[0], gpcOutL2_22[1], gpcOutL2_21[2]}, gpcOutL3_29);
gpc015 gpcL3_30 ({gpcOutL2_133[0], gpcOutL2_115[2], gpcOutL2_91[0], gpcOutL2_25[0], gpcOutL2_24[1], gpcOutL2_23[2]}, gpcOutL3_30);
gpc015 gpcL3_31 ({gpcOutL2_117[1], gpcOutL2_117[0], gpcOutL2_116[2], gpcOutL2_52[0], gpcOutL2_51[1], gpcOutL2_50[2]}, gpcOutL3_31);
gpc015 gpcL3_32 ({gpcOutL2_118[1], gpcOutL2_118[0], gpcOutL2_117[2], gpcOutL2_54[0], gpcOutL2_53[1], gpcOutL2_52[2]}, gpcOutL3_32);
gpc015 gpcL3_33 ({gpcOutL2_119[1], gpcOutL2_119[0], gpcOutL2_118[2], gpcOutL2_56[0], gpcOutL2_55[1], gpcOutL2_54[2]}, gpcOutL3_33);
gpc015 gpcL3_34 ({gpcOutL2_120[1], gpcOutL2_120[0], gpcOutL2_119[2], gpcOutL2_58[0], gpcOutL2_57[1], gpcOutL2_56[2]}, gpcOutL3_34);
gpc015 gpcL3_35 ({gpcOutL2_127[1], gpcOutL2_127[0], gpcOutL2_120[2], gpcOutL2_60[0], gpcOutL2_59[1], gpcOutL2_58[2]}, gpcOutL3_35);
gpc015 gpcL3_36 ({gpcOutL2_139[0], gpcOutL2_127[3], gpcOutL2_63[0], gpcOutL2_62[1], gpcOutL2_61[2], gpcOutL1_75[2]}, gpcOutL3_36);
gpc015 gpcL3_37 ({gpcOutL2_67[0], gpcOutL2_139[2], gpcOutL2_66[0], gpcOutL2_65[1], gpcOutL2_64[2], pp255[5]}, gpcOutL3_37);
gpc005 gpcL3_38 ({gpcOutL2_93[1], gpcOutL2_76[0], gpcOutL2_30[0], gpcOutL2_29[1], gpcOutL2_28[2]}, gpcOutL3_38);
gpc005 gpcL3_39 ({gpcOutL2_136[0], gpcOutL2_95[1], gpcOutL2_47[0], gpcOutL2_46[1], gpcOutL2_45[2]}, gpcOutL3_39);
gpc005 gpcL3_40 ({gpcOutL2_110[0], gpcOutL2_96[1], gpcOutL2_49[0], gpcOutL2_48[1], gpcOutL2_47[2]}, gpcOutL3_40);
gpc014 gpcL3_41 ({gpcOutL2_113[2], gpcOutL2_113[1], gpcOutL2_106[2], gpcOutL1_5[1], gpcOutL1_4[2]}, gpcOutL3_41);
gpc014 gpcL3_42 ({gpcOutL2_5[0], gpcOutL2_101[2], gpcOutL2_4[0], gpcOutL2_3[1], pp7[5]}, gpcOutL3_42);
gpc014 gpcL3_43 ({gpcOutL2_7[0], gpcOutL2_6[0], gpcOutL2_5[1], gpcOutL2_4[2], gpcOutL0_25[2]}, gpcOutL3_43);
gpc014 gpcL3_44 ({gpcOutL2_126[1], gpcOutL2_126[0], gpcOutL2_11[0], gpcOutL2_10[1], gpcOutL2_9[2]}, gpcOutL3_44);
gpc014 gpcL3_45 ({gpcOutL2_137[1], gpcOutL2_137[0], gpcOutL2_97[1], gpcOutL2_75[2], gpcOutL0_96[2]}, gpcOutL3_45);
gpc023 gpcL3_46 ({gpcOutL2_8[0], gpcOutL2_7[1], gpcOutL2_6[1], gpcOutL2_5[2], gpcOutL1_19[2]}, gpcOutL3_46);
gpc023 gpcL3_47 ({gpcOutL2_126[2], gpcOutL2_13[0], gpcOutL2_12[0], gpcOutL2_11[1], gpcOutL2_10[2]}, gpcOutL3_47);
gpc023 gpcL3_48 ({gpcOutL2_127[2], gpcOutL2_62[0], gpcOutL2_61[0], gpcOutL2_60[1], gpcOutL2_59[2]}, gpcOutL3_48);
gpc023 gpcL3_49 ({gpcOutL2_139[1], gpcOutL2_65[0], gpcOutL2_64[0], gpcOutL2_63[1], gpcOutL2_62[2]}, gpcOutL3_49);
gpc023 gpcL3_50 ({gpcOutL2_69[0], gpcOutL2_68[1], gpcOutL2_68[0], gpcOutL2_67[1], gpcOutL2_66[2]}, gpcOutL3_50);
gpc023 gpcL3_51 ({gpcOutL2_71[0], gpcOutL2_70[1], gpcOutL2_70[0], gpcOutL2_69[1], gpcOutL2_68[2]}, gpcOutL3_51);
gpc023 gpcL3_52 ({gpcOutL2_73[0], gpcOutL2_72[1], gpcOutL2_72[0], gpcOutL2_71[1], gpcOutL2_70[2]}, gpcOutL3_52);
gpc023 gpcL3_53 ({gpcOutL2_75[0], gpcOutL2_74[1], gpcOutL2_74[0], gpcOutL2_73[1], gpcOutL2_72[2]}, gpcOutL3_53);
gpc003 gpcL3_54 ({gpcOutL2_4[1], gpcOutL2_3[2], gpcOutL0_24[2]}, gpcOutL3_54);
gpc003 gpcL3_55 ({gpcOutL2_9[1], gpcOutL2_8[2], gpcOutL1_22[2]}, gpcOutL3_55);
gpc003 gpcL3_56 ({gpcOutL2_15[0], gpcOutL2_14[1], gpcOutL2_13[2]}, gpcOutL3_56);
gpc003 gpcL3_57 ({gpcOutL2_17[0], gpcOutL2_16[1], gpcOutL2_15[2]}, gpcOutL3_57);
gpc003 gpcL3_58 ({gpcOutL2_131[0], gpcOutL2_19[0], gpcOutL2_18[1]}, gpcOutL3_58);
gpc003 gpcL3_59 ({gpcOutL2_108[1], gpcOutL2_21[0], gpcOutL2_20[1]}, gpcOutL3_59);
gpc003 gpcL3_60 ({gpcOutL2_91[1], gpcOutL2_26[0], gpcOutL2_25[1]}, gpcOutL3_60);
gpc003 gpcL3_61 ({gpcOutL2_53[0], gpcOutL2_52[1], gpcOutL2_51[2]}, gpcOutL3_61);
gpc003 gpcL3_62 ({gpcOutL2_55[0], gpcOutL2_54[1], gpcOutL2_53[2]}, gpcOutL3_62);
gpc003 gpcL3_63 ({gpcOutL2_57[0], gpcOutL2_56[1], gpcOutL2_55[2]}, gpcOutL3_63);
gpc003 gpcL3_64 ({gpcOutL2_59[0], gpcOutL2_58[1], gpcOutL2_57[2]}, gpcOutL3_64);
gpc003 gpcL3_65 ({gpcOutL2_97[0], gpcOutL2_75[1], gpcOutL2_74[2]}, gpcOutL3_65);
gpc023 gpcL3_66 ({gpcOutL2_140[3], gpcOutL1_228[0], gpcOutL2_140[2], gpcOutL0_448[2], gpcOutL0_0[0]}, gpcOutL3_66);

// level 4
wire [2:0]  gpcOutL4_0;
wire [2:0]  gpcOutL4_1;
wire [2:0]  gpcOutL4_2;
wire [2:0]  gpcOutL4_3;
wire [2:0]  gpcOutL4_4;
wire [2:0]  gpcOutL4_5;
wire [2:0]  gpcOutL4_6;
wire [2:0]  gpcOutL4_7;
wire [2:0]  gpcOutL4_8;
wire [2:0]  gpcOutL4_9;
wire [2:0]  gpcOutL4_10;
wire [2:0]  gpcOutL4_11;
wire [2:0]  gpcOutL4_12;
wire [2:0]  gpcOutL4_13;
wire [2:0]  gpcOutL4_14;
wire [2:0]  gpcOutL4_15;
wire [2:0]  gpcOutL4_16;
wire [2:0]  gpcOutL4_17;
wire [3:0]  gpcOutL4_18;

gpc014 gpcL4_0 ({gpcOutL3_46[2], gpcOutL3_46[1], gpcOutL3_43[2], gpcOutL2_6[2], gpcOutL1_20[2]}, gpcOutL4_0);
gpc014 gpcL4_1 ({gpcOutL3_47[2], gpcOutL3_47[1], gpcOutL3_44[2], gpcOutL2_12[1], gpcOutL2_11[2]}, gpcOutL4_1);
gpc014 gpcL4_2 ({gpcOutL3_60[1], gpcOutL3_60[0], gpcOutL3_30[1], gpcOutL3_2[2], gpcOutL2_24[2]}, gpcOutL4_2);
gpc014 gpcL4_3 ({gpcOutL3_21[0], gpcOutL3_20[0], gpcOutL3_19[1], gpcOutL3_18[2], gpcOutL0_64[2]}, gpcOutL4_3);
gpc014 gpcL4_4 ({gpcOutL3_61[1], gpcOutL3_61[0], gpcOutL3_31[1], gpcOutL3_24[2], gpcOutL1_65[2]}, gpcOutL4_4);
gpc014 gpcL4_5 ({gpcOutL3_48[2], gpcOutL3_48[1], gpcOutL3_35[2], gpcOutL2_61[1], gpcOutL2_60[2]}, gpcOutL4_5);
gpc014 gpcL4_6 ({gpcOutL3_49[2], gpcOutL3_49[1], gpcOutL3_36[2], gpcOutL2_64[1], gpcOutL2_63[2]}, gpcOutL4_6);
gpc023 gpcL4_7 ({gpcOutL3_56[1], gpcOutL3_27[0], gpcOutL3_56[0], gpcOutL3_26[1], gpcOutL1_27[2]}, gpcOutL4_7);
gpc023 gpcL4_8 ({gpcOutL3_57[1], gpcOutL3_27[2], gpcOutL3_57[0], gpcOutL3_27[1], gpcOutL1_29[2]}, gpcOutL4_8);
gpc023 gpcL4_9 ({gpcOutL3_58[1], gpcOutL3_28[0], gpcOutL3_58[0], gpcOutL3_0[1], gpcOutL2_17[2]}, gpcOutL4_9);
gpc023 gpcL4_10 ({gpcOutL3_59[1], gpcOutL3_28[2], gpcOutL3_59[0], gpcOutL3_28[1], gpcOutL2_19[2]}, gpcOutL4_10);
gpc023 gpcL4_11 ({gpcOutL3_39[1], gpcOutL3_22[0], gpcOutL3_39[0], gpcOutL3_21[1], gpcOutL3_20[2]}, gpcOutL4_11);
gpc023 gpcL4_12 ({gpcOutL3_40[1], gpcOutL3_23[0], gpcOutL3_40[0], gpcOutL3_39[2], gpcOutL3_22[1]}, gpcOutL4_12);
gpc023 gpcL4_13 ({gpcOutL3_31[0], gpcOutL3_24[1], gpcOutL3_40[2], gpcOutL3_24[0], gpcOutL3_23[1]}, gpcOutL4_13);
gpc023 gpcL4_14 ({gpcOutL3_62[1], gpcOutL3_33[0], gpcOutL3_62[0], gpcOutL3_32[1], gpcOutL1_67[2]}, gpcOutL4_14);
gpc023 gpcL4_15 ({gpcOutL3_63[1], gpcOutL3_34[0], gpcOutL3_63[0], gpcOutL3_33[1], gpcOutL1_69[2]}, gpcOutL4_15);
gpc023 gpcL4_16 ({gpcOutL3_64[1], gpcOutL3_35[0], gpcOutL3_64[0], gpcOutL3_34[1], gpcOutL0_78[2]}, gpcOutL4_16);
gpc023 gpcL4_17 ({gpcOutL3_50[0], gpcOutL3_37[2], gpcOutL3_37[1], gpcOutL2_66[1], gpcOutL2_65[2]}, gpcOutL4_17);
gpc213 gpcL4_18 ({gpcOutL2_104[1], gpcOutL1_216[0], gpcOutL2_104[0], gpcOutL3_66[2], gpcOutL1_236[0], gpcOutL1_228[1]}, gpcOutL4_18);

// final adder
wire [114:0]  adderIn0;
wire [114:0]  adderIn1;
wire [114:0]  adderIn2;
wire [115:0]  adderOut;

assign adderIn0 = {pp511[5], gpcOutL1_265[1], gpcOutL1_265[0], gpcOutL1_254[1], gpcOutL1_254[0], gpcOutL1_253[1], gpcOutL2_125[2], gpcOutL2_125[1], gpcOutL2_125[0], gpcOutL2_124[1], gpcOutL2_124[0], gpcOutL2_123[1], gpcOutL2_123[0], gpcOutL2_122[1], gpcOutL2_122[0], gpcOutL2_121[1], gpcOutL2_121[0], gpcOutL2_111[0], gpcOutL2_138[1], gpcOutL3_45[2], gpcOutL3_45[1], gpcOutL3_65[1], gpcOutL3_65[0], gpcOutL3_53[1], gpcOutL3_53[0], gpcOutL3_52[1], gpcOutL3_52[0], gpcOutL3_51[1], gpcOutL3_51[0], gpcOutL4_17[2], gpcOutL4_17[1], gpcOutL4_17[0], gpcOutL4_6[1], gpcOutL4_6[0], gpcOutL4_5[2], gpcOutL4_5[1], gpcOutL4_5[0], gpcOutL4_16[2], gpcOutL4_16[1], gpcOutL4_16[0], gpcOutL4_15[1], gpcOutL4_15[0], gpcOutL4_14[1], gpcOutL4_14[0], gpcOutL4_4[1], gpcOutL4_13[2], gpcOutL4_13[1], gpcOutL4_13[0], gpcOutL4_12[1], gpcOutL4_12[0], gpcOutL4_11[1], gpcOutL4_11[0], gpcOutL4_3[1], gpcOutL4_3[0], gpcOutL3_19[0], gpcOutL3_18[0], gpcOutL3_17[0], gpcOutL3_16[0], gpcOutL3_15[0], gpcOutL3_14[0], gpcOutL3_13[0], gpcOutL3_12[0], gpcOutL3_11[0], gpcOutL3_10[0], gpcOutL3_9[0], gpcOutL3_8[0], gpcOutL3_38[2], gpcOutL3_38[1], gpcOutL3_38[0], gpcOutL3_5[0], gpcOutL4_2[2], gpcOutL4_2[1], gpcOutL4_2[0], gpcOutL3_30[0], gpcOutL3_29[1], gpcOutL4_10[2], gpcOutL4_10[1], gpcOutL4_10[0], gpcOutL4_9[1], gpcOutL4_9[0], gpcOutL4_8[1], gpcOutL4_8[0], gpcOutL4_7[1], gpcOutL4_7[0], gpcOutL4_1[1], gpcOutL4_1[0], gpcOutL3_47[0], gpcOutL3_55[1], gpcOutL4_0[2], gpcOutL4_0[1], gpcOutL4_0[0], gpcOutL3_46[0], gpcOutL3_54[1], gpcOutL3_54[0], gpcOutL3_42[0], gpcOutL2_101[1], gpcOutL2_101[0], gpcOutL2_100[2], gpcOutL2_100[1], gpcOutL2_100[0], gpcOutL2_90[1], gpcOutL2_130[1], gpcOutL2_130[0], gpcOutL2_129[1], gpcOutL3_41[2], gpcOutL3_41[1], gpcOutL3_41[0], gpcOutL2_113[0], gpcOutL2_128[1], gpcOutL2_128[0], gpcOutL2_105[0], gpcOutL1_220[1], gpcOutL2_112[2], gpcOutL2_112[1], gpcOutL4_18[3]};
assign adderIn1 = {1'b0, pp511[4], gpcOutL1_254[2], 1'b0, gpcOutL1_253[2], gpcOutL0_463[2], gpcOutL1_253[0], gpcOutL0_110[2], gpcOutL2_124[2], gpcOutL1_101[1], gpcOutL2_123[2], gpcOutL1_99[2], gpcOutL2_122[2], gpcOutL1_97[2], gpcOutL2_121[2], gpcOutL2_111[2], gpcOutL2_111[1], gpcOutL2_99[1], gpcOutL2_99[0], gpcOutL2_138[0], gpcOutL2_98[0], gpcOutL3_45[0], gpcOutL3_53[2], gpcOutL2_73[2], gpcOutL3_52[2], gpcOutL2_71[2], gpcOutL3_51[2], gpcOutL2_69[2], gpcOutL3_50[2], gpcOutL3_50[1], 1'b0, gpcOutL4_6[2], gpcOutL3_37[0], 1'b0, gpcOutL3_49[0], gpcOutL3_36[0], 1'b0, gpcOutL3_48[0], gpcOutL3_34[2], gpcOutL4_15[2], gpcOutL3_33[2], gpcOutL4_14[2], gpcOutL3_32[2], gpcOutL4_4[2], gpcOutL3_32[0], gpcOutL4_4[0], gpcOutL3_23[2], gpcOutL4_12[2], gpcOutL3_22[2], gpcOutL4_11[2], gpcOutL3_21[2], gpcOutL4_3[2], gpcOutL3_20[1], 1'b0, gpcOutL3_18[1], gpcOutL3_17[1], gpcOutL3_16[1], gpcOutL3_15[1], gpcOutL3_14[1], gpcOutL3_13[1], gpcOutL3_12[1], gpcOutL3_11[1], gpcOutL3_10[1], gpcOutL3_9[1], gpcOutL3_8[1], gpcOutL3_7[1], gpcOutL3_7[0], gpcOutL3_6[0], gpcOutL3_5[1], gpcOutL3_4[1], gpcOutL3_4[0], gpcOutL3_30[2], 1'b0, gpcOutL3_29[2], gpcOutL3_2[0], gpcOutL3_29[0], gpcOutL3_1[0], gpcOutL4_9[2], gpcOutL3_0[2], gpcOutL4_8[2], gpcOutL3_0[0], gpcOutL4_7[2], gpcOutL3_26[2], gpcOutL4_1[2], gpcOutL3_26[0], 1'b0, gpcOutL3_44[1], gpcOutL3_44[0], gpcOutL3_55[0], gpcOutL3_25[0], 1'b0, gpcOutL3_43[1], gpcOutL3_43[0], gpcOutL3_42[1], 1'b0, gpcOutL2_3[0], gpcOutL2_2[1], gpcOutL2_2[0], gpcOutL2_1[0], gpcOutL2_90[2], gpcOutL2_0[0], gpcOutL2_90[0], gpcOutL2_89[1], gpcOutL2_89[0], gpcOutL2_129[0], gpcOutL2_88[0], 1'b0, gpcOutL2_106[1], gpcOutL2_106[0], gpcOutL2_105[1], 1'b0, gpcOutL1_1[0], gpcOutL1_220[0], gpcOutL1_0[0], gpcOutL2_112[0]};
assign adderIn2 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, gpcOutL1_252[2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, gpcOutL1_95[2], gpcOutL2_99[2], 1'b0, gpcOutL2_98[2], gpcOutL2_98[1], gpcOutL2_97[2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, gpcOutL2_67[2], 1'b0, 1'b0, 1'b0, 1'b0, gpcOutL3_36[1], 1'b0, 1'b0, gpcOutL3_35[1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, gpcOutL3_31[2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, gpcOutL3_19[2], 1'b0, gpcOutL3_17[2], gpcOutL3_16[2], gpcOutL3_15[2], gpcOutL3_14[2], gpcOutL3_13[2], gpcOutL3_12[2], gpcOutL3_11[2], gpcOutL3_10[2], gpcOutL3_9[2], gpcOutL3_8[2], gpcOutL3_7[2], gpcOutL3_6[2], gpcOutL3_6[1], gpcOutL3_5[2], gpcOutL3_4[2], gpcOutL3_3[2], gpcOutL3_3[1], gpcOutL3_3[0], 1'b0, gpcOutL3_2[1], gpcOutL3_1[2], gpcOutL3_1[1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, gpcOutL3_25[2], gpcOutL3_25[1], 1'b0, 1'b0, 1'b0, gpcOutL3_42[2], 1'b0, 1'b0, gpcOutL2_2[2], gpcOutL2_1[2], gpcOutL2_1[1], gpcOutL2_0[2], gpcOutL2_0[1], 1'b0, gpcOutL2_89[2], gpcOutL1_8[2], gpcOutL2_88[2], gpcOutL2_88[1], 1'b0, 1'b0, 1'b0, gpcOutL2_105[2], 1'b0, 1'b0, gpcOutL1_0[2], gpcOutL1_0[1], 1'b0, gpcOutL2_104[2]};
assign adderOut = adderIn0 + adderIn1 + adderIn2;

// multiplayer output
assign out = {adderOut[114:0], gpcOutL4_18[2], gpcOutL4_18[1], gpcOutL4_18[0], gpcOutL3_66[1], gpcOutL3_66[0], gpcOutL2_140[1], gpcOutL2_140[0], gpcOutL1_269[1], gpcOutL1_269[0], gpcOutL0_519[1], gpcOutL0_519[0], pp0[1], pp0[0]};

endmodule


/******************************************/

