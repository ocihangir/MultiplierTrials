module mult_32x64_lut6_akak(in0, in1, out);

input  [31:0]  in0;
input  [63:0]  in1;
output  [95:0]  out;

wire [5:0]  pp0;
wire [5:0]  pp1;
wire [5:0]  pp2;
wire [5:0]  pp3;
wire [5:0]  pp4;
wire [5:0]  pp5;
wire [5:0]  pp6;
wire [5:0]  pp7;
wire [5:0]  pp8;
wire [5:0]  pp9;
wire [5:0]  pp10;
wire [5:0]  pp11;
wire [5:0]  pp12;
wire [5:0]  pp13;
wire [5:0]  pp14;
wire [5:0]  pp15;
wire [5:0]  pp16;
wire [5:0]  pp17;
wire [5:0]  pp18;
wire [5:0]  pp19;
wire [5:0]  pp20;
wire [5:0]  pp21;
wire [5:0]  pp22;
wire [5:0]  pp23;
wire [5:0]  pp24;
wire [5:0]  pp25;
wire [5:0]  pp26;
wire [5:0]  pp27;
wire [5:0]  pp28;
wire [5:0]  pp29;
wire [5:0]  pp30;
wire [5:0]  pp31;
wire [5:0]  pp32;
wire [5:0]  pp33;
wire [5:0]  pp34;
wire [5:0]  pp35;
wire [5:0]  pp36;
wire [5:0]  pp37;
wire [5:0]  pp38;
wire [5:0]  pp39;
wire [5:0]  pp40;
wire [5:0]  pp41;
wire [5:0]  pp42;
wire [5:0]  pp43;
wire [5:0]  pp44;
wire [5:0]  pp45;
wire [5:0]  pp46;
wire [5:0]  pp47;
wire [5:0]  pp48;
wire [5:0]  pp49;
wire [5:0]  pp50;
wire [5:0]  pp51;
wire [5:0]  pp52;
wire [5:0]  pp53;
wire [5:0]  pp54;
wire [5:0]  pp55;
wire [5:0]  pp56;
wire [5:0]  pp57;
wire [5:0]  pp58;
wire [5:0]  pp59;
wire [5:0]  pp60;
wire [5:0]  pp61;
wire [5:0]  pp62;
wire [5:0]  pp63;
wire [5:0]  pp64;
wire [5:0]  pp65;
wire [5:0]  pp66;
wire [5:0]  pp67;
wire [5:0]  pp68;
wire [5:0]  pp69;
wire [5:0]  pp70;
wire [5:0]  pp71;
wire [5:0]  pp72;
wire [5:0]  pp73;
wire [5:0]  pp74;
wire [5:0]  pp75;
wire [5:0]  pp76;
wire [5:0]  pp77;
wire [5:0]  pp78;
wire [5:0]  pp79;
wire [5:0]  pp80;
wire [5:0]  pp81;
wire [5:0]  pp82;
wire [5:0]  pp83;
wire [5:0]  pp84;
wire [5:0]  pp85;
wire [5:0]  pp86;
wire [5:0]  pp87;
wire [5:0]  pp88;
wire [5:0]  pp89;
wire [5:0]  pp90;
wire [5:0]  pp91;
wire [5:0]  pp92;
wire [5:0]  pp93;
wire [5:0]  pp94;
wire [5:0]  pp95;
wire [5:0]  pp96;
wire [5:0]  pp97;
wire [5:0]  pp98;
wire [5:0]  pp99;
wire [5:0]  pp100;
wire [5:0]  pp101;
wire [5:0]  pp102;
wire [5:0]  pp103;
wire [5:0]  pp104;
wire [5:0]  pp105;
wire [5:0]  pp106;
wire [5:0]  pp107;
wire [5:0]  pp108;
wire [5:0]  pp109;
wire [5:0]  pp110;
wire [5:0]  pp111;
wire [5:0]  pp112;
wire [5:0]  pp113;
wire [5:0]  pp114;
wire [5:0]  pp115;
wire [5:0]  pp116;
wire [5:0]  pp117;
wire [5:0]  pp118;
wire [5:0]  pp119;
wire [5:0]  pp120;
wire [5:0]  pp121;
wire [5:0]  pp122;
wire [5:0]  pp123;
wire [5:0]  pp124;
wire [5:0]  pp125;
wire [5:0]  pp126;
wire [5:0]  pp127;
wire [5:0]  pp128;
wire [5:0]  pp129;
wire [5:0]  pp130;
wire [5:0]  pp131;
wire [5:0]  pp132;
wire [5:0]  pp133;
wire [5:0]  pp134;
wire [5:0]  pp135;
wire [5:0]  pp136;
wire [5:0]  pp137;
wire [5:0]  pp138;
wire [5:0]  pp139;
wire [5:0]  pp140;
wire [5:0]  pp141;
wire [5:0]  pp142;
wire [5:0]  pp143;
wire [5:0]  pp144;
wire [5:0]  pp145;
wire [5:0]  pp146;
wire [5:0]  pp147;
wire [5:0]  pp148;
wire [5:0]  pp149;
wire [5:0]  pp150;
wire [5:0]  pp151;
wire [5:0]  pp152;
wire [5:0]  pp153;
wire [5:0]  pp154;
wire [5:0]  pp155;
wire [5:0]  pp156;
wire [5:0]  pp157;
wire [5:0]  pp158;
wire [5:0]  pp159;
wire [5:0]  pp160;
wire [5:0]  pp161;
wire [5:0]  pp162;
wire [5:0]  pp163;
wire [5:0]  pp164;
wire [5:0]  pp165;
wire [5:0]  pp166;
wire [5:0]  pp167;
wire [5:0]  pp168;
wire [5:0]  pp169;
wire [5:0]  pp170;
wire [5:0]  pp171;
wire [5:0]  pp172;
wire [5:0]  pp173;
wire [5:0]  pp174;
wire [5:0]  pp175;
wire [5:0]  pp176;
wire [5:0]  pp177;
wire [5:0]  pp178;
wire [5:0]  pp179;
wire [5:0]  pp180;
wire [5:0]  pp181;
wire [5:0]  pp182;
wire [5:0]  pp183;
wire [5:0]  pp184;
wire [5:0]  pp185;
wire [5:0]  pp186;
wire [5:0]  pp187;
wire [5:0]  pp188;
wire [5:0]  pp189;
wire [5:0]  pp190;
wire [5:0]  pp191;
wire [5:0]  pp192;
wire [5:0]  pp193;
wire [5:0]  pp194;
wire [5:0]  pp195;
wire [5:0]  pp196;
wire [5:0]  pp197;
wire [5:0]  pp198;
wire [5:0]  pp199;
wire [5:0]  pp200;
wire [5:0]  pp201;
wire [5:0]  pp202;
wire [5:0]  pp203;
wire [5:0]  pp204;
wire [5:0]  pp205;
wire [5:0]  pp206;
wire [5:0]  pp207;
wire [5:0]  pp208;
wire [5:0]  pp209;
wire [5:0]  pp210;
wire [5:0]  pp211;
wire [5:0]  pp212;
wire [5:0]  pp213;
wire [5:0]  pp214;
wire [5:0]  pp215;
wire [5:0]  pp216;
wire [5:0]  pp217;
wire [5:0]  pp218;
wire [5:0]  pp219;
wire [5:0]  pp220;
wire [5:0]  pp221;
wire [5:0]  pp222;
wire [5:0]  pp223;
wire [5:0]  pp224;
wire [5:0]  pp225;
wire [5:0]  pp226;
wire [5:0]  pp227;
wire [5:0]  pp228;
wire [5:0]  pp229;
wire [5:0]  pp230;
wire [5:0]  pp231;
wire [5:0]  pp232;
wire [5:0]  pp233;
wire [5:0]  pp234;
wire [5:0]  pp235;
wire [5:0]  pp236;
wire [5:0]  pp237;
wire [5:0]  pp238;
wire [5:0]  pp239;
wire [5:0]  pp240;
wire [5:0]  pp241;
wire [5:0]  pp242;
wire [5:0]  pp243;
wire [5:0]  pp244;
wire [5:0]  pp245;
wire [5:0]  pp246;
wire [5:0]  pp247;
wire [5:0]  pp248;
wire [5:0]  pp249;
wire [5:0]  pp250;
wire [5:0]  pp251;
wire [5:0]  pp252;
wire [5:0]  pp253;
wire [5:0]  pp254;
wire [5:0]  pp255;

// partial products
level0_mult lvl0_mult0({in0[3:0], in1[1:0]}, pp0);
level0_mult lvl0_mult1({in0[7:4], in1[1:0]}, pp1);
level0_mult lvl0_mult2({in0[11:8], in1[1:0]}, pp2);
level0_mult lvl0_mult3({in0[15:12], in1[1:0]}, pp3);
level0_mult lvl0_mult4({in0[19:16], in1[1:0]}, pp4);
level0_mult lvl0_mult5({in0[23:20], in1[1:0]}, pp5);
level0_mult lvl0_mult6({in0[27:24], in1[1:0]}, pp6);
level0_mult lvl0_mult7({in0[31:28], in1[1:0]}, pp7);
level0_mult lvl0_mult8({in0[3:0], in1[3:2]}, pp8);
level0_mult lvl0_mult9({in0[7:4], in1[3:2]}, pp9);
level0_mult lvl0_mult10({in0[11:8], in1[3:2]}, pp10);
level0_mult lvl0_mult11({in0[15:12], in1[3:2]}, pp11);
level0_mult lvl0_mult12({in0[19:16], in1[3:2]}, pp12);
level0_mult lvl0_mult13({in0[23:20], in1[3:2]}, pp13);
level0_mult lvl0_mult14({in0[27:24], in1[3:2]}, pp14);
level0_mult lvl0_mult15({in0[31:28], in1[3:2]}, pp15);
level0_mult lvl0_mult16({in0[3:0], in1[5:4]}, pp16);
level0_mult lvl0_mult17({in0[7:4], in1[5:4]}, pp17);
level0_mult lvl0_mult18({in0[11:8], in1[5:4]}, pp18);
level0_mult lvl0_mult19({in0[15:12], in1[5:4]}, pp19);
level0_mult lvl0_mult20({in0[19:16], in1[5:4]}, pp20);
level0_mult lvl0_mult21({in0[23:20], in1[5:4]}, pp21);
level0_mult lvl0_mult22({in0[27:24], in1[5:4]}, pp22);
level0_mult lvl0_mult23({in0[31:28], in1[5:4]}, pp23);
level0_mult lvl0_mult24({in0[3:0], in1[7:6]}, pp24);
level0_mult lvl0_mult25({in0[7:4], in1[7:6]}, pp25);
level0_mult lvl0_mult26({in0[11:8], in1[7:6]}, pp26);
level0_mult lvl0_mult27({in0[15:12], in1[7:6]}, pp27);
level0_mult lvl0_mult28({in0[19:16], in1[7:6]}, pp28);
level0_mult lvl0_mult29({in0[23:20], in1[7:6]}, pp29);
level0_mult lvl0_mult30({in0[27:24], in1[7:6]}, pp30);
level0_mult lvl0_mult31({in0[31:28], in1[7:6]}, pp31);
level0_mult lvl0_mult32({in0[3:0], in1[9:8]}, pp32);
level0_mult lvl0_mult33({in0[7:4], in1[9:8]}, pp33);
level0_mult lvl0_mult34({in0[11:8], in1[9:8]}, pp34);
level0_mult lvl0_mult35({in0[15:12], in1[9:8]}, pp35);
level0_mult lvl0_mult36({in0[19:16], in1[9:8]}, pp36);
level0_mult lvl0_mult37({in0[23:20], in1[9:8]}, pp37);
level0_mult lvl0_mult38({in0[27:24], in1[9:8]}, pp38);
level0_mult lvl0_mult39({in0[31:28], in1[9:8]}, pp39);
level0_mult lvl0_mult40({in0[3:0], in1[11:10]}, pp40);
level0_mult lvl0_mult41({in0[7:4], in1[11:10]}, pp41);
level0_mult lvl0_mult42({in0[11:8], in1[11:10]}, pp42);
level0_mult lvl0_mult43({in0[15:12], in1[11:10]}, pp43);
level0_mult lvl0_mult44({in0[19:16], in1[11:10]}, pp44);
level0_mult lvl0_mult45({in0[23:20], in1[11:10]}, pp45);
level0_mult lvl0_mult46({in0[27:24], in1[11:10]}, pp46);
level0_mult lvl0_mult47({in0[31:28], in1[11:10]}, pp47);
level0_mult lvl0_mult48({in0[3:0], in1[13:12]}, pp48);
level0_mult lvl0_mult49({in0[7:4], in1[13:12]}, pp49);
level0_mult lvl0_mult50({in0[11:8], in1[13:12]}, pp50);
level0_mult lvl0_mult51({in0[15:12], in1[13:12]}, pp51);
level0_mult lvl0_mult52({in0[19:16], in1[13:12]}, pp52);
level0_mult lvl0_mult53({in0[23:20], in1[13:12]}, pp53);
level0_mult lvl0_mult54({in0[27:24], in1[13:12]}, pp54);
level0_mult lvl0_mult55({in0[31:28], in1[13:12]}, pp55);
level0_mult lvl0_mult56({in0[3:0], in1[15:14]}, pp56);
level0_mult lvl0_mult57({in0[7:4], in1[15:14]}, pp57);
level0_mult lvl0_mult58({in0[11:8], in1[15:14]}, pp58);
level0_mult lvl0_mult59({in0[15:12], in1[15:14]}, pp59);
level0_mult lvl0_mult60({in0[19:16], in1[15:14]}, pp60);
level0_mult lvl0_mult61({in0[23:20], in1[15:14]}, pp61);
level0_mult lvl0_mult62({in0[27:24], in1[15:14]}, pp62);
level0_mult lvl0_mult63({in0[31:28], in1[15:14]}, pp63);
level0_mult lvl0_mult64({in0[3:0], in1[17:16]}, pp64);
level0_mult lvl0_mult65({in0[7:4], in1[17:16]}, pp65);
level0_mult lvl0_mult66({in0[11:8], in1[17:16]}, pp66);
level0_mult lvl0_mult67({in0[15:12], in1[17:16]}, pp67);
level0_mult lvl0_mult68({in0[19:16], in1[17:16]}, pp68);
level0_mult lvl0_mult69({in0[23:20], in1[17:16]}, pp69);
level0_mult lvl0_mult70({in0[27:24], in1[17:16]}, pp70);
level0_mult lvl0_mult71({in0[31:28], in1[17:16]}, pp71);
level0_mult lvl0_mult72({in0[3:0], in1[19:18]}, pp72);
level0_mult lvl0_mult73({in0[7:4], in1[19:18]}, pp73);
level0_mult lvl0_mult74({in0[11:8], in1[19:18]}, pp74);
level0_mult lvl0_mult75({in0[15:12], in1[19:18]}, pp75);
level0_mult lvl0_mult76({in0[19:16], in1[19:18]}, pp76);
level0_mult lvl0_mult77({in0[23:20], in1[19:18]}, pp77);
level0_mult lvl0_mult78({in0[27:24], in1[19:18]}, pp78);
level0_mult lvl0_mult79({in0[31:28], in1[19:18]}, pp79);
level0_mult lvl0_mult80({in0[3:0], in1[21:20]}, pp80);
level0_mult lvl0_mult81({in0[7:4], in1[21:20]}, pp81);
level0_mult lvl0_mult82({in0[11:8], in1[21:20]}, pp82);
level0_mult lvl0_mult83({in0[15:12], in1[21:20]}, pp83);
level0_mult lvl0_mult84({in0[19:16], in1[21:20]}, pp84);
level0_mult lvl0_mult85({in0[23:20], in1[21:20]}, pp85);
level0_mult lvl0_mult86({in0[27:24], in1[21:20]}, pp86);
level0_mult lvl0_mult87({in0[31:28], in1[21:20]}, pp87);
level0_mult lvl0_mult88({in0[3:0], in1[23:22]}, pp88);
level0_mult lvl0_mult89({in0[7:4], in1[23:22]}, pp89);
level0_mult lvl0_mult90({in0[11:8], in1[23:22]}, pp90);
level0_mult lvl0_mult91({in0[15:12], in1[23:22]}, pp91);
level0_mult lvl0_mult92({in0[19:16], in1[23:22]}, pp92);
level0_mult lvl0_mult93({in0[23:20], in1[23:22]}, pp93);
level0_mult lvl0_mult94({in0[27:24], in1[23:22]}, pp94);
level0_mult lvl0_mult95({in0[31:28], in1[23:22]}, pp95);
level0_mult lvl0_mult96({in0[3:0], in1[25:24]}, pp96);
level0_mult lvl0_mult97({in0[7:4], in1[25:24]}, pp97);
level0_mult lvl0_mult98({in0[11:8], in1[25:24]}, pp98);
level0_mult lvl0_mult99({in0[15:12], in1[25:24]}, pp99);
level0_mult lvl0_mult100({in0[19:16], in1[25:24]}, pp100);
level0_mult lvl0_mult101({in0[23:20], in1[25:24]}, pp101);
level0_mult lvl0_mult102({in0[27:24], in1[25:24]}, pp102);
level0_mult lvl0_mult103({in0[31:28], in1[25:24]}, pp103);
level0_mult lvl0_mult104({in0[3:0], in1[27:26]}, pp104);
level0_mult lvl0_mult105({in0[7:4], in1[27:26]}, pp105);
level0_mult lvl0_mult106({in0[11:8], in1[27:26]}, pp106);
level0_mult lvl0_mult107({in0[15:12], in1[27:26]}, pp107);
level0_mult lvl0_mult108({in0[19:16], in1[27:26]}, pp108);
level0_mult lvl0_mult109({in0[23:20], in1[27:26]}, pp109);
level0_mult lvl0_mult110({in0[27:24], in1[27:26]}, pp110);
level0_mult lvl0_mult111({in0[31:28], in1[27:26]}, pp111);
level0_mult lvl0_mult112({in0[3:0], in1[29:28]}, pp112);
level0_mult lvl0_mult113({in0[7:4], in1[29:28]}, pp113);
level0_mult lvl0_mult114({in0[11:8], in1[29:28]}, pp114);
level0_mult lvl0_mult115({in0[15:12], in1[29:28]}, pp115);
level0_mult lvl0_mult116({in0[19:16], in1[29:28]}, pp116);
level0_mult lvl0_mult117({in0[23:20], in1[29:28]}, pp117);
level0_mult lvl0_mult118({in0[27:24], in1[29:28]}, pp118);
level0_mult lvl0_mult119({in0[31:28], in1[29:28]}, pp119);
level0_mult lvl0_mult120({in0[3:0], in1[31:30]}, pp120);
level0_mult lvl0_mult121({in0[7:4], in1[31:30]}, pp121);
level0_mult lvl0_mult122({in0[11:8], in1[31:30]}, pp122);
level0_mult lvl0_mult123({in0[15:12], in1[31:30]}, pp123);
level0_mult lvl0_mult124({in0[19:16], in1[31:30]}, pp124);
level0_mult lvl0_mult125({in0[23:20], in1[31:30]}, pp125);
level0_mult lvl0_mult126({in0[27:24], in1[31:30]}, pp126);
level0_mult lvl0_mult127({in0[31:28], in1[31:30]}, pp127);
level0_mult lvl0_mult128({in0[3:0], in1[33:32]}, pp128);
level0_mult lvl0_mult129({in0[7:4], in1[33:32]}, pp129);
level0_mult lvl0_mult130({in0[11:8], in1[33:32]}, pp130);
level0_mult lvl0_mult131({in0[15:12], in1[33:32]}, pp131);
level0_mult lvl0_mult132({in0[19:16], in1[33:32]}, pp132);
level0_mult lvl0_mult133({in0[23:20], in1[33:32]}, pp133);
level0_mult lvl0_mult134({in0[27:24], in1[33:32]}, pp134);
level0_mult lvl0_mult135({in0[31:28], in1[33:32]}, pp135);
level0_mult lvl0_mult136({in0[3:0], in1[35:34]}, pp136);
level0_mult lvl0_mult137({in0[7:4], in1[35:34]}, pp137);
level0_mult lvl0_mult138({in0[11:8], in1[35:34]}, pp138);
level0_mult lvl0_mult139({in0[15:12], in1[35:34]}, pp139);
level0_mult lvl0_mult140({in0[19:16], in1[35:34]}, pp140);
level0_mult lvl0_mult141({in0[23:20], in1[35:34]}, pp141);
level0_mult lvl0_mult142({in0[27:24], in1[35:34]}, pp142);
level0_mult lvl0_mult143({in0[31:28], in1[35:34]}, pp143);
level0_mult lvl0_mult144({in0[3:0], in1[37:36]}, pp144);
level0_mult lvl0_mult145({in0[7:4], in1[37:36]}, pp145);
level0_mult lvl0_mult146({in0[11:8], in1[37:36]}, pp146);
level0_mult lvl0_mult147({in0[15:12], in1[37:36]}, pp147);
level0_mult lvl0_mult148({in0[19:16], in1[37:36]}, pp148);
level0_mult lvl0_mult149({in0[23:20], in1[37:36]}, pp149);
level0_mult lvl0_mult150({in0[27:24], in1[37:36]}, pp150);
level0_mult lvl0_mult151({in0[31:28], in1[37:36]}, pp151);
level0_mult lvl0_mult152({in0[3:0], in1[39:38]}, pp152);
level0_mult lvl0_mult153({in0[7:4], in1[39:38]}, pp153);
level0_mult lvl0_mult154({in0[11:8], in1[39:38]}, pp154);
level0_mult lvl0_mult155({in0[15:12], in1[39:38]}, pp155);
level0_mult lvl0_mult156({in0[19:16], in1[39:38]}, pp156);
level0_mult lvl0_mult157({in0[23:20], in1[39:38]}, pp157);
level0_mult lvl0_mult158({in0[27:24], in1[39:38]}, pp158);
level0_mult lvl0_mult159({in0[31:28], in1[39:38]}, pp159);
level0_mult lvl0_mult160({in0[3:0], in1[41:40]}, pp160);
level0_mult lvl0_mult161({in0[7:4], in1[41:40]}, pp161);
level0_mult lvl0_mult162({in0[11:8], in1[41:40]}, pp162);
level0_mult lvl0_mult163({in0[15:12], in1[41:40]}, pp163);
level0_mult lvl0_mult164({in0[19:16], in1[41:40]}, pp164);
level0_mult lvl0_mult165({in0[23:20], in1[41:40]}, pp165);
level0_mult lvl0_mult166({in0[27:24], in1[41:40]}, pp166);
level0_mult lvl0_mult167({in0[31:28], in1[41:40]}, pp167);
level0_mult lvl0_mult168({in0[3:0], in1[43:42]}, pp168);
level0_mult lvl0_mult169({in0[7:4], in1[43:42]}, pp169);
level0_mult lvl0_mult170({in0[11:8], in1[43:42]}, pp170);
level0_mult lvl0_mult171({in0[15:12], in1[43:42]}, pp171);
level0_mult lvl0_mult172({in0[19:16], in1[43:42]}, pp172);
level0_mult lvl0_mult173({in0[23:20], in1[43:42]}, pp173);
level0_mult lvl0_mult174({in0[27:24], in1[43:42]}, pp174);
level0_mult lvl0_mult175({in0[31:28], in1[43:42]}, pp175);
level0_mult lvl0_mult176({in0[3:0], in1[45:44]}, pp176);
level0_mult lvl0_mult177({in0[7:4], in1[45:44]}, pp177);
level0_mult lvl0_mult178({in0[11:8], in1[45:44]}, pp178);
level0_mult lvl0_mult179({in0[15:12], in1[45:44]}, pp179);
level0_mult lvl0_mult180({in0[19:16], in1[45:44]}, pp180);
level0_mult lvl0_mult181({in0[23:20], in1[45:44]}, pp181);
level0_mult lvl0_mult182({in0[27:24], in1[45:44]}, pp182);
level0_mult lvl0_mult183({in0[31:28], in1[45:44]}, pp183);
level0_mult lvl0_mult184({in0[3:0], in1[47:46]}, pp184);
level0_mult lvl0_mult185({in0[7:4], in1[47:46]}, pp185);
level0_mult lvl0_mult186({in0[11:8], in1[47:46]}, pp186);
level0_mult lvl0_mult187({in0[15:12], in1[47:46]}, pp187);
level0_mult lvl0_mult188({in0[19:16], in1[47:46]}, pp188);
level0_mult lvl0_mult189({in0[23:20], in1[47:46]}, pp189);
level0_mult lvl0_mult190({in0[27:24], in1[47:46]}, pp190);
level0_mult lvl0_mult191({in0[31:28], in1[47:46]}, pp191);
level0_mult lvl0_mult192({in0[3:0], in1[49:48]}, pp192);
level0_mult lvl0_mult193({in0[7:4], in1[49:48]}, pp193);
level0_mult lvl0_mult194({in0[11:8], in1[49:48]}, pp194);
level0_mult lvl0_mult195({in0[15:12], in1[49:48]}, pp195);
level0_mult lvl0_mult196({in0[19:16], in1[49:48]}, pp196);
level0_mult lvl0_mult197({in0[23:20], in1[49:48]}, pp197);
level0_mult lvl0_mult198({in0[27:24], in1[49:48]}, pp198);
level0_mult lvl0_mult199({in0[31:28], in1[49:48]}, pp199);
level0_mult lvl0_mult200({in0[3:0], in1[51:50]}, pp200);
level0_mult lvl0_mult201({in0[7:4], in1[51:50]}, pp201);
level0_mult lvl0_mult202({in0[11:8], in1[51:50]}, pp202);
level0_mult lvl0_mult203({in0[15:12], in1[51:50]}, pp203);
level0_mult lvl0_mult204({in0[19:16], in1[51:50]}, pp204);
level0_mult lvl0_mult205({in0[23:20], in1[51:50]}, pp205);
level0_mult lvl0_mult206({in0[27:24], in1[51:50]}, pp206);
level0_mult lvl0_mult207({in0[31:28], in1[51:50]}, pp207);
level0_mult lvl0_mult208({in0[3:0], in1[53:52]}, pp208);
level0_mult lvl0_mult209({in0[7:4], in1[53:52]}, pp209);
level0_mult lvl0_mult210({in0[11:8], in1[53:52]}, pp210);
level0_mult lvl0_mult211({in0[15:12], in1[53:52]}, pp211);
level0_mult lvl0_mult212({in0[19:16], in1[53:52]}, pp212);
level0_mult lvl0_mult213({in0[23:20], in1[53:52]}, pp213);
level0_mult lvl0_mult214({in0[27:24], in1[53:52]}, pp214);
level0_mult lvl0_mult215({in0[31:28], in1[53:52]}, pp215);
level0_mult lvl0_mult216({in0[3:0], in1[55:54]}, pp216);
level0_mult lvl0_mult217({in0[7:4], in1[55:54]}, pp217);
level0_mult lvl0_mult218({in0[11:8], in1[55:54]}, pp218);
level0_mult lvl0_mult219({in0[15:12], in1[55:54]}, pp219);
level0_mult lvl0_mult220({in0[19:16], in1[55:54]}, pp220);
level0_mult lvl0_mult221({in0[23:20], in1[55:54]}, pp221);
level0_mult lvl0_mult222({in0[27:24], in1[55:54]}, pp222);
level0_mult lvl0_mult223({in0[31:28], in1[55:54]}, pp223);
level0_mult lvl0_mult224({in0[3:0], in1[57:56]}, pp224);
level0_mult lvl0_mult225({in0[7:4], in1[57:56]}, pp225);
level0_mult lvl0_mult226({in0[11:8], in1[57:56]}, pp226);
level0_mult lvl0_mult227({in0[15:12], in1[57:56]}, pp227);
level0_mult lvl0_mult228({in0[19:16], in1[57:56]}, pp228);
level0_mult lvl0_mult229({in0[23:20], in1[57:56]}, pp229);
level0_mult lvl0_mult230({in0[27:24], in1[57:56]}, pp230);
level0_mult lvl0_mult231({in0[31:28], in1[57:56]}, pp231);
level0_mult lvl0_mult232({in0[3:0], in1[59:58]}, pp232);
level0_mult lvl0_mult233({in0[7:4], in1[59:58]}, pp233);
level0_mult lvl0_mult234({in0[11:8], in1[59:58]}, pp234);
level0_mult lvl0_mult235({in0[15:12], in1[59:58]}, pp235);
level0_mult lvl0_mult236({in0[19:16], in1[59:58]}, pp236);
level0_mult lvl0_mult237({in0[23:20], in1[59:58]}, pp237);
level0_mult lvl0_mult238({in0[27:24], in1[59:58]}, pp238);
level0_mult lvl0_mult239({in0[31:28], in1[59:58]}, pp239);
level0_mult lvl0_mult240({in0[3:0], in1[61:60]}, pp240);
level0_mult lvl0_mult241({in0[7:4], in1[61:60]}, pp241);
level0_mult lvl0_mult242({in0[11:8], in1[61:60]}, pp242);
level0_mult lvl0_mult243({in0[15:12], in1[61:60]}, pp243);
level0_mult lvl0_mult244({in0[19:16], in1[61:60]}, pp244);
level0_mult lvl0_mult245({in0[23:20], in1[61:60]}, pp245);
level0_mult lvl0_mult246({in0[27:24], in1[61:60]}, pp246);
level0_mult lvl0_mult247({in0[31:28], in1[61:60]}, pp247);
level0_mult lvl0_mult248({in0[3:0], in1[63:62]}, pp248);
level0_mult lvl0_mult249({in0[7:4], in1[63:62]}, pp249);
level0_mult lvl0_mult250({in0[11:8], in1[63:62]}, pp250);
level0_mult lvl0_mult251({in0[15:12], in1[63:62]}, pp251);
level0_mult lvl0_mult252({in0[19:16], in1[63:62]}, pp252);
level0_mult lvl0_mult253({in0[23:20], in1[63:62]}, pp253);
level0_mult lvl0_mult254({in0[27:24], in1[63:62]}, pp254);
level0_mult lvl0_mult255({in0[31:28], in1[63:62]}, pp255);


// level 0
wire [2:0]  gpcOutL0_0;
wire [2:0]  gpcOutL0_1;
wire [2:0]  gpcOutL0_2;
wire [2:0]  gpcOutL0_3;
wire [2:0]  gpcOutL0_4;
wire [2:0]  gpcOutL0_5;
wire [2:0]  gpcOutL0_6;
wire [2:0]  gpcOutL0_7;
wire [2:0]  gpcOutL0_8;
wire [2:0]  gpcOutL0_9;
wire [2:0]  gpcOutL0_10;
wire [2:0]  gpcOutL0_11;
wire [2:0]  gpcOutL0_12;
wire [2:0]  gpcOutL0_13;
wire [2:0]  gpcOutL0_14;
wire [2:0]  gpcOutL0_15;
wire [2:0]  gpcOutL0_16;
wire [2:0]  gpcOutL0_17;
wire [2:0]  gpcOutL0_18;
wire [2:0]  gpcOutL0_19;
wire [2:0]  gpcOutL0_20;
wire [2:0]  gpcOutL0_21;
wire [2:0]  gpcOutL0_22;
wire [2:0]  gpcOutL0_23;
wire [2:0]  gpcOutL0_24;
wire [2:0]  gpcOutL0_25;
wire [2:0]  gpcOutL0_26;
wire [2:0]  gpcOutL0_27;
wire [2:0]  gpcOutL0_28;
wire [2:0]  gpcOutL0_29;
wire [2:0]  gpcOutL0_30;
wire [2:0]  gpcOutL0_31;
wire [2:0]  gpcOutL0_32;
wire [2:0]  gpcOutL0_33;
wire [2:0]  gpcOutL0_34;
wire [2:0]  gpcOutL0_35;
wire [2:0]  gpcOutL0_36;
wire [2:0]  gpcOutL0_37;
wire [2:0]  gpcOutL0_38;
wire [2:0]  gpcOutL0_39;
wire [2:0]  gpcOutL0_40;
wire [2:0]  gpcOutL0_41;
wire [2:0]  gpcOutL0_42;
wire [2:0]  gpcOutL0_43;
wire [2:0]  gpcOutL0_44;
wire [2:0]  gpcOutL0_45;
wire [2:0]  gpcOutL0_46;
wire [2:0]  gpcOutL0_47;
wire [2:0]  gpcOutL0_48;
wire [2:0]  gpcOutL0_49;
wire [2:0]  gpcOutL0_50;
wire [2:0]  gpcOutL0_51;
wire [2:0]  gpcOutL0_52;
wire [2:0]  gpcOutL0_53;
wire [2:0]  gpcOutL0_54;
wire [2:0]  gpcOutL0_55;
wire [2:0]  gpcOutL0_56;
wire [2:0]  gpcOutL0_57;
wire [2:0]  gpcOutL0_58;
wire [2:0]  gpcOutL0_59;
wire [2:0]  gpcOutL0_60;
wire [2:0]  gpcOutL0_61;
wire [2:0]  gpcOutL0_62;
wire [2:0]  gpcOutL0_63;
wire [2:0]  gpcOutL0_64;
wire [2:0]  gpcOutL0_65;
wire [2:0]  gpcOutL0_66;
wire [2:0]  gpcOutL0_67;
wire [2:0]  gpcOutL0_68;
wire [2:0]  gpcOutL0_69;
wire [2:0]  gpcOutL0_70;
wire [2:0]  gpcOutL0_71;
wire [2:0]  gpcOutL0_72;
wire [2:0]  gpcOutL0_73;
wire [2:0]  gpcOutL0_74;
wire [2:0]  gpcOutL0_75;
wire [2:0]  gpcOutL0_76;
wire [2:0]  gpcOutL0_77;
wire [2:0]  gpcOutL0_78;
wire [2:0]  gpcOutL0_79;
wire [2:0]  gpcOutL0_80;
wire [2:0]  gpcOutL0_81;
wire [2:0]  gpcOutL0_82;
wire [2:0]  gpcOutL0_83;
wire [2:0]  gpcOutL0_84;
wire [2:0]  gpcOutL0_85;
wire [2:0]  gpcOutL0_86;
wire [2:0]  gpcOutL0_87;
wire [2:0]  gpcOutL0_88;
wire [2:0]  gpcOutL0_89;
wire [2:0]  gpcOutL0_90;
wire [2:0]  gpcOutL0_91;
wire [2:0]  gpcOutL0_92;
wire [2:0]  gpcOutL0_93;
wire [2:0]  gpcOutL0_94;
wire [2:0]  gpcOutL0_95;
wire [2:0]  gpcOutL0_96;
wire [2:0]  gpcOutL0_97;
wire [2:0]  gpcOutL0_98;
wire [2:0]  gpcOutL0_99;
wire [2:0]  gpcOutL0_100;
wire [2:0]  gpcOutL0_101;
wire [2:0]  gpcOutL0_102;
wire [2:0]  gpcOutL0_103;
wire [2:0]  gpcOutL0_104;
wire [2:0]  gpcOutL0_105;
wire [2:0]  gpcOutL0_106;
wire [2:0]  gpcOutL0_107;
wire [2:0]  gpcOutL0_108;
wire [2:0]  gpcOutL0_109;
wire [2:0]  gpcOutL0_110;
wire [2:0]  gpcOutL0_111;
wire [2:0]  gpcOutL0_112;
wire [2:0]  gpcOutL0_113;
wire [2:0]  gpcOutL0_114;
wire [2:0]  gpcOutL0_115;
wire [2:0]  gpcOutL0_116;
wire [2:0]  gpcOutL0_117;
wire [2:0]  gpcOutL0_118;
wire [2:0]  gpcOutL0_119;
wire [2:0]  gpcOutL0_120;
wire [2:0]  gpcOutL0_121;
wire [2:0]  gpcOutL0_122;
wire [2:0]  gpcOutL0_123;
wire [2:0]  gpcOutL0_124;
wire [2:0]  gpcOutL0_125;
wire [2:0]  gpcOutL0_126;
wire [2:0]  gpcOutL0_127;
wire [2:0]  gpcOutL0_128;
wire [2:0]  gpcOutL0_129;
wire [2:0]  gpcOutL0_130;
wire [2:0]  gpcOutL0_131;
wire [2:0]  gpcOutL0_132;
wire [2:0]  gpcOutL0_133;
wire [2:0]  gpcOutL0_134;
wire [2:0]  gpcOutL0_135;
wire [2:0]  gpcOutL0_136;
wire [2:0]  gpcOutL0_137;
wire [2:0]  gpcOutL0_138;
wire [2:0]  gpcOutL0_139;
wire [2:0]  gpcOutL0_140;
wire [2:0]  gpcOutL0_141;
wire [2:0]  gpcOutL0_142;
wire [2:0]  gpcOutL0_143;
wire [2:0]  gpcOutL0_144;
wire [2:0]  gpcOutL0_145;
wire [2:0]  gpcOutL0_146;
wire [2:0]  gpcOutL0_147;
wire [2:0]  gpcOutL0_148;
wire [2:0]  gpcOutL0_149;
wire [2:0]  gpcOutL0_150;
wire [2:0]  gpcOutL0_151;
wire [2:0]  gpcOutL0_152;
wire [2:0]  gpcOutL0_153;
wire [2:0]  gpcOutL0_154;
wire [2:0]  gpcOutL0_155;
wire [2:0]  gpcOutL0_156;
wire [2:0]  gpcOutL0_157;
wire [2:0]  gpcOutL0_158;
wire [2:0]  gpcOutL0_159;
wire [2:0]  gpcOutL0_160;
wire [2:0]  gpcOutL0_161;
wire [2:0]  gpcOutL0_162;
wire [2:0]  gpcOutL0_163;
wire [2:0]  gpcOutL0_164;
wire [2:0]  gpcOutL0_165;
wire [2:0]  gpcOutL0_166;
wire [2:0]  gpcOutL0_167;
wire [2:0]  gpcOutL0_168;
wire [2:0]  gpcOutL0_169;
wire [2:0]  gpcOutL0_170;
wire [2:0]  gpcOutL0_171;
wire [2:0]  gpcOutL0_172;
wire [2:0]  gpcOutL0_173;
wire [2:0]  gpcOutL0_174;
wire [2:0]  gpcOutL0_175;
wire [2:0]  gpcOutL0_176;
wire [2:0]  gpcOutL0_177;
wire [2:0]  gpcOutL0_178;
wire [2:0]  gpcOutL0_179;
wire [2:0]  gpcOutL0_180;
wire [2:0]  gpcOutL0_181;
wire [2:0]  gpcOutL0_182;
wire [2:0]  gpcOutL0_183;
wire [2:0]  gpcOutL0_184;
wire [2:0]  gpcOutL0_185;
wire [2:0]  gpcOutL0_186;
wire [2:0]  gpcOutL0_187;
wire [2:0]  gpcOutL0_188;
wire [2:0]  gpcOutL0_189;
wire [2:0]  gpcOutL0_190;
wire [2:0]  gpcOutL0_191;
wire [2:0]  gpcOutL0_192;
wire [2:0]  gpcOutL0_193;
wire [2:0]  gpcOutL0_194;
wire [2:0]  gpcOutL0_195;
wire [2:0]  gpcOutL0_196;
wire [2:0]  gpcOutL0_197;
wire [2:0]  gpcOutL0_198;
wire [2:0]  gpcOutL0_199;
wire [2:0]  gpcOutL0_200;
wire [2:0]  gpcOutL0_201;
wire [2:0]  gpcOutL0_202;
wire [2:0]  gpcOutL0_203;
wire [2:0]  gpcOutL0_204;
wire [2:0]  gpcOutL0_205;
wire [2:0]  gpcOutL0_206;
wire [2:0]  gpcOutL0_207;
wire [2:0]  gpcOutL0_208;
wire [2:0]  gpcOutL0_209;
wire [2:0]  gpcOutL0_210;
wire [2:0]  gpcOutL0_211;
wire [2:0]  gpcOutL0_212;
wire [2:0]  gpcOutL0_213;
wire [2:0]  gpcOutL0_214;
wire [2:0]  gpcOutL0_215;
wire [2:0]  gpcOutL0_216;
wire [2:0]  gpcOutL0_217;
wire [2:0]  gpcOutL0_218;
wire [2:0]  gpcOutL0_219;
wire [2:0]  gpcOutL0_220;
wire [2:0]  gpcOutL0_221;
wire [2:0]  gpcOutL0_222;
wire [2:0]  gpcOutL0_223;
wire [2:0]  gpcOutL0_224;
wire [2:0]  gpcOutL0_225;
wire [2:0]  gpcOutL0_226;
wire [2:0]  gpcOutL0_227;
wire [2:0]  gpcOutL0_228;
wire [2:0]  gpcOutL0_229;
wire [2:0]  gpcOutL0_230;
wire [2:0]  gpcOutL0_231;
wire [2:0]  gpcOutL0_232;
wire [2:0]  gpcOutL0_233;
wire [2:0]  gpcOutL0_234;
wire [2:0]  gpcOutL0_235;
wire [2:0]  gpcOutL0_236;
wire [2:0]  gpcOutL0_237;
wire [2:0]  gpcOutL0_238;
wire [2:0]  gpcOutL0_239;
wire [2:0]  gpcOutL0_240;
wire [2:0]  gpcOutL0_241;
wire [2:0]  gpcOutL0_242;
wire [2:0]  gpcOutL0_243;
wire [2:0]  gpcOutL0_244;
wire [2:0]  gpcOutL0_245;
wire [2:0]  gpcOutL0_246;
wire [1:0]  gpcOutL0_247;
wire [1:0]  gpcOutL0_248;
wire [1:0]  gpcOutL0_249;
wire [1:0]  gpcOutL0_250;
wire [1:0]  gpcOutL0_251;
wire [1:0]  gpcOutL0_252;
wire [1:0]  gpcOutL0_253;
wire [1:0]  gpcOutL0_254;
wire [1:0]  gpcOutL0_255;
wire [2:0]  gpcOutL0_256;
wire [2:0]  gpcOutL0_257;
wire [2:0]  gpcOutL0_258;
wire [2:0]  gpcOutL0_259;

gpc006 gpcL0_0 ({pp32[0], pp24[2], pp17[0], pp16[4], pp9[2], pp2[0]}, gpcOutL0_0);
gpc006 gpcL0_1 ({pp32[1], pp24[3], pp17[1], pp16[5], pp9[3], pp2[1]}, gpcOutL0_1);
gpc006 gpcL0_2 ({pp40[0], pp32[2], pp25[0], pp24[4], pp17[2], pp10[0]}, gpcOutL0_2);
gpc006 gpcL0_3 ({pp40[1], pp32[3], pp25[1], pp24[5], pp17[3], pp10[1]}, gpcOutL0_3);
gpc006 gpcL0_4 ({pp48[0], pp40[2], pp33[0], pp32[4], pp25[2], pp18[0]}, gpcOutL0_4);
gpc006 gpcL0_5 ({pp48[1], pp40[3], pp33[1], pp32[5], pp25[3], pp18[1]}, gpcOutL0_5);
gpc006 gpcL0_6 ({pp56[0], pp48[2], pp41[0], pp40[4], pp33[2], pp26[0]}, gpcOutL0_6);
gpc006 gpcL0_7 ({pp56[1], pp48[3], pp41[1], pp40[5], pp33[3], pp26[1]}, gpcOutL0_7);
gpc006 gpcL0_8 ({pp64[0], pp56[2], pp49[0], pp48[4], pp41[2], pp34[0]}, gpcOutL0_8);
gpc006 gpcL0_9 ({pp64[1], pp56[3], pp49[1], pp48[5], pp41[3], pp34[1]}, gpcOutL0_9);
gpc006 gpcL0_10 ({pp72[0], pp64[2], pp57[0], pp56[4], pp49[2], pp42[0]}, gpcOutL0_10);
gpc006 gpcL0_11 ({pp72[1], pp64[3], pp57[1], pp56[5], pp49[3], pp42[1]}, gpcOutL0_11);
gpc006 gpcL0_12 ({pp80[0], pp72[2], pp65[0], pp64[4], pp57[2], pp50[0]}, gpcOutL0_12);
gpc006 gpcL0_13 ({pp80[1], pp72[3], pp65[1], pp64[5], pp57[3], pp50[1]}, gpcOutL0_13);
gpc006 gpcL0_14 ({pp88[0], pp80[2], pp73[0], pp72[4], pp65[2], pp58[0]}, gpcOutL0_14);
gpc006 gpcL0_15 ({pp88[1], pp80[3], pp73[1], pp72[5], pp65[3], pp58[1]}, gpcOutL0_15);
gpc006 gpcL0_16 ({pp96[0], pp88[2], pp81[0], pp80[4], pp73[2], pp66[0]}, gpcOutL0_16);
gpc006 gpcL0_17 ({pp96[1], pp88[3], pp81[1], pp80[5], pp73[3], pp66[1]}, gpcOutL0_17);
gpc006 gpcL0_18 ({pp104[0], pp96[2], pp89[0], pp88[4], pp81[2], pp74[0]}, gpcOutL0_18);
gpc006 gpcL0_19 ({pp104[1], pp96[3], pp89[1], pp88[5], pp81[3], pp74[1]}, gpcOutL0_19);
gpc006 gpcL0_20 ({pp112[0], pp104[2], pp97[0], pp96[4], pp89[2], pp82[0]}, gpcOutL0_20);
gpc006 gpcL0_21 ({pp112[1], pp104[3], pp97[1], pp96[5], pp89[3], pp82[1]}, gpcOutL0_21);
gpc006 gpcL0_22 ({pp120[0], pp112[2], pp105[0], pp104[4], pp97[2], pp90[0]}, gpcOutL0_22);
gpc006 gpcL0_23 ({pp120[1], pp112[3], pp105[1], pp104[5], pp97[3], pp90[1]}, gpcOutL0_23);
gpc006 gpcL0_24 ({pp128[0], pp120[2], pp113[0], pp112[4], pp105[2], pp98[0]}, gpcOutL0_24);
gpc006 gpcL0_25 ({pp128[1], pp120[3], pp113[1], pp112[5], pp105[3], pp98[1]}, gpcOutL0_25);
gpc006 gpcL0_26 ({pp136[0], pp128[2], pp121[0], pp120[4], pp113[2], pp106[0]}, gpcOutL0_26);
gpc006 gpcL0_27 ({pp136[1], pp128[3], pp121[1], pp120[5], pp113[3], pp106[1]}, gpcOutL0_27);
gpc006 gpcL0_28 ({pp144[0], pp136[2], pp129[0], pp128[4], pp121[2], pp114[0]}, gpcOutL0_28);
gpc006 gpcL0_29 ({pp144[1], pp136[3], pp129[1], pp128[5], pp121[3], pp114[1]}, gpcOutL0_29);
gpc006 gpcL0_30 ({pp152[0], pp144[2], pp137[0], pp136[4], pp129[2], pp122[0]}, gpcOutL0_30);
gpc006 gpcL0_31 ({pp152[1], pp144[3], pp137[1], pp136[5], pp129[3], pp122[1]}, gpcOutL0_31);
gpc006 gpcL0_32 ({pp160[0], pp152[2], pp145[0], pp144[4], pp137[2], pp130[0]}, gpcOutL0_32);
gpc006 gpcL0_33 ({pp160[1], pp152[3], pp145[1], pp144[5], pp137[3], pp130[1]}, gpcOutL0_33);
gpc006 gpcL0_34 ({pp168[0], pp160[2], pp153[0], pp152[4], pp145[2], pp138[0]}, gpcOutL0_34);
gpc006 gpcL0_35 ({pp168[1], pp160[3], pp153[1], pp152[5], pp145[3], pp138[1]}, gpcOutL0_35);
gpc006 gpcL0_36 ({pp176[0], pp168[2], pp161[0], pp160[4], pp153[2], pp146[0]}, gpcOutL0_36);
gpc006 gpcL0_37 ({pp176[1], pp168[3], pp161[1], pp160[5], pp153[3], pp146[1]}, gpcOutL0_37);
gpc006 gpcL0_38 ({pp184[0], pp176[2], pp169[0], pp168[4], pp161[2], pp154[0]}, gpcOutL0_38);
gpc006 gpcL0_39 ({pp184[1], pp176[3], pp169[1], pp168[5], pp161[3], pp154[1]}, gpcOutL0_39);
gpc006 gpcL0_40 ({pp192[0], pp184[2], pp177[0], pp176[4], pp169[2], pp162[0]}, gpcOutL0_40);
gpc006 gpcL0_41 ({pp192[1], pp184[3], pp177[1], pp176[5], pp169[3], pp162[1]}, gpcOutL0_41);
gpc006 gpcL0_42 ({pp200[0], pp192[2], pp185[0], pp184[4], pp177[2], pp170[0]}, gpcOutL0_42);
gpc006 gpcL0_43 ({pp200[1], pp192[3], pp185[1], pp184[5], pp177[3], pp170[1]}, gpcOutL0_43);
gpc006 gpcL0_44 ({pp208[0], pp200[2], pp193[0], pp192[4], pp185[2], pp178[0]}, gpcOutL0_44);
gpc006 gpcL0_45 ({pp208[1], pp200[3], pp193[1], pp192[5], pp185[3], pp178[1]}, gpcOutL0_45);
gpc006 gpcL0_46 ({pp216[0], pp208[2], pp201[0], pp200[4], pp193[2], pp186[0]}, gpcOutL0_46);
gpc006 gpcL0_47 ({pp216[1], pp208[3], pp201[1], pp200[5], pp193[3], pp186[1]}, gpcOutL0_47);
gpc006 gpcL0_48 ({pp224[0], pp216[2], pp209[0], pp208[4], pp201[2], pp194[0]}, gpcOutL0_48);
gpc006 gpcL0_49 ({pp224[1], pp216[3], pp209[1], pp208[5], pp201[3], pp194[1]}, gpcOutL0_49);
gpc006 gpcL0_50 ({pp232[0], pp224[2], pp217[0], pp216[4], pp209[2], pp202[0]}, gpcOutL0_50);
gpc006 gpcL0_51 ({pp232[1], pp224[3], pp217[1], pp216[5], pp209[3], pp202[1]}, gpcOutL0_51);
gpc006 gpcL0_52 ({pp240[0], pp232[2], pp225[0], pp224[4], pp217[2], pp210[0]}, gpcOutL0_52);
gpc006 gpcL0_53 ({pp240[1], pp232[3], pp225[1], pp224[5], pp217[3], pp210[1]}, gpcOutL0_53);
gpc006 gpcL0_54 ({pp248[0], pp240[2], pp233[0], pp232[4], pp225[2], pp218[0]}, gpcOutL0_54);
gpc006 gpcL0_55 ({pp248[1], pp240[3], pp233[1], pp232[5], pp225[3], pp218[1]}, gpcOutL0_55);
gpc006 gpcL0_56 ({pp248[2], pp241[0], pp240[4], pp233[2], pp226[0], pp225[4]}, gpcOutL0_56);
gpc006 gpcL0_57 ({pp248[3], pp241[1], pp240[5], pp233[3], pp226[1], pp225[5]}, gpcOutL0_57);
gpc006 gpcL0_58 ({pp249[0], pp248[4], pp241[2], pp234[0], pp233[4], pp226[2]}, gpcOutL0_58);
gpc006 gpcL0_59 ({pp249[1], pp248[5], pp241[3], pp234[1], pp233[5], pp226[3]}, gpcOutL0_59);
gpc006 gpcL0_60 ({pp249[2], pp242[0], pp241[4], pp234[2], pp227[0], pp226[4]}, gpcOutL0_60);
gpc006 gpcL0_61 ({pp249[3], pp242[1], pp241[5], pp234[3], pp227[1], pp226[5]}, gpcOutL0_61);
gpc006 gpcL0_62 ({pp250[0], pp249[4], pp242[2], pp235[0], pp234[4], pp227[2]}, gpcOutL0_62);
gpc006 gpcL0_63 ({pp250[1], pp249[5], pp242[3], pp235[1], pp234[5], pp227[3]}, gpcOutL0_63);
gpc006 gpcL0_64 ({pp250[2], pp243[0], pp242[4], pp235[2], pp228[0], pp227[4]}, gpcOutL0_64);
gpc006 gpcL0_65 ({pp250[3], pp243[1], pp242[5], pp235[3], pp228[1], pp227[5]}, gpcOutL0_65);
gpc006 gpcL0_66 ({pp251[0], pp250[4], pp243[2], pp236[0], pp235[4], pp228[2]}, gpcOutL0_66);
gpc006 gpcL0_67 ({pp251[1], pp250[5], pp243[3], pp236[1], pp235[5], pp228[3]}, gpcOutL0_67);
gpc006 gpcL0_68 ({pp251[2], pp244[0], pp243[4], pp236[2], pp229[0], pp228[4]}, gpcOutL0_68);
gpc006 gpcL0_69 ({pp251[3], pp244[1], pp243[5], pp236[3], pp229[1], pp228[5]}, gpcOutL0_69);
gpc006 gpcL0_70 ({pp252[0], pp251[4], pp244[2], pp237[0], pp236[4], pp229[2]}, gpcOutL0_70);
gpc006 gpcL0_71 ({pp252[1], pp251[5], pp244[3], pp237[1], pp236[5], pp229[3]}, gpcOutL0_71);
gpc006 gpcL0_72 ({pp252[2], pp245[0], pp244[4], pp237[2], pp230[0], pp229[4]}, gpcOutL0_72);
gpc006 gpcL0_73 ({pp252[3], pp245[1], pp244[5], pp237[3], pp230[1], pp229[5]}, gpcOutL0_73);
gpc006 gpcL0_74 ({pp253[0], pp252[4], pp245[2], pp238[0], pp237[4], pp230[2]}, gpcOutL0_74);
gpc006 gpcL0_75 ({pp253[1], pp252[5], pp245[3], pp238[1], pp237[5], pp230[3]}, gpcOutL0_75);
gpc006 gpcL0_76 ({pp253[2], pp246[0], pp245[4], pp238[2], pp231[0], pp230[4]}, gpcOutL0_76);
gpc006 gpcL0_77 ({pp253[3], pp246[1], pp245[5], pp238[3], pp231[1], pp230[5]}, gpcOutL0_77);
gpc006 gpcL0_78 ({pp254[0], pp253[4], pp246[2], pp239[0], pp238[4], pp231[2]}, gpcOutL0_78);
gpc006 gpcL0_79 ({pp254[1], pp253[5], pp246[3], pp239[1], pp238[5], pp231[3]}, gpcOutL0_79);
gpc006 gpcL0_80 ({pp33[4], pp26[2], pp19[0], pp18[4], pp11[2], pp4[0]}, gpcOutL0_80);
gpc006 gpcL0_81 ({pp33[5], pp26[3], pp19[1], pp18[5], pp11[3], pp4[1]}, gpcOutL0_81);
gpc006 gpcL0_82 ({pp41[4], pp34[2], pp27[0], pp26[4], pp19[2], pp12[0]}, gpcOutL0_82);
gpc006 gpcL0_83 ({pp41[5], pp34[3], pp27[1], pp26[5], pp19[3], pp12[1]}, gpcOutL0_83);
gpc006 gpcL0_84 ({pp49[4], pp42[2], pp35[0], pp34[4], pp27[2], pp20[0]}, gpcOutL0_84);
gpc006 gpcL0_85 ({pp49[5], pp42[3], pp35[1], pp34[5], pp27[3], pp20[1]}, gpcOutL0_85);
gpc006 gpcL0_86 ({pp57[4], pp50[2], pp43[0], pp42[4], pp35[2], pp28[0]}, gpcOutL0_86);
gpc006 gpcL0_87 ({pp57[5], pp50[3], pp43[1], pp42[5], pp35[3], pp28[1]}, gpcOutL0_87);
gpc006 gpcL0_88 ({pp65[4], pp58[2], pp51[0], pp50[4], pp43[2], pp36[0]}, gpcOutL0_88);
gpc006 gpcL0_89 ({pp65[5], pp58[3], pp51[1], pp50[5], pp43[3], pp36[1]}, gpcOutL0_89);
gpc006 gpcL0_90 ({pp73[4], pp66[2], pp59[0], pp58[4], pp51[2], pp44[0]}, gpcOutL0_90);
gpc006 gpcL0_91 ({pp73[5], pp66[3], pp59[1], pp58[5], pp51[3], pp44[1]}, gpcOutL0_91);
gpc006 gpcL0_92 ({pp81[4], pp74[2], pp67[0], pp66[4], pp59[2], pp52[0]}, gpcOutL0_92);
gpc006 gpcL0_93 ({pp81[5], pp74[3], pp67[1], pp66[5], pp59[3], pp52[1]}, gpcOutL0_93);
gpc006 gpcL0_94 ({pp89[4], pp82[2], pp75[0], pp74[4], pp67[2], pp60[0]}, gpcOutL0_94);
gpc006 gpcL0_95 ({pp89[5], pp82[3], pp75[1], pp74[5], pp67[3], pp60[1]}, gpcOutL0_95);
gpc006 gpcL0_96 ({pp97[4], pp90[2], pp83[0], pp82[4], pp75[2], pp68[0]}, gpcOutL0_96);
gpc006 gpcL0_97 ({pp97[5], pp90[3], pp83[1], pp82[5], pp75[3], pp68[1]}, gpcOutL0_97);
gpc006 gpcL0_98 ({pp105[4], pp98[2], pp91[0], pp90[4], pp83[2], pp76[0]}, gpcOutL0_98);
gpc006 gpcL0_99 ({pp105[5], pp98[3], pp91[1], pp90[5], pp83[3], pp76[1]}, gpcOutL0_99);
gpc006 gpcL0_100 ({pp113[4], pp106[2], pp99[0], pp98[4], pp91[2], pp84[0]}, gpcOutL0_100);
gpc006 gpcL0_101 ({pp113[5], pp106[3], pp99[1], pp98[5], pp91[3], pp84[1]}, gpcOutL0_101);
gpc006 gpcL0_102 ({pp121[4], pp114[2], pp107[0], pp106[4], pp99[2], pp92[0]}, gpcOutL0_102);
gpc006 gpcL0_103 ({pp121[5], pp114[3], pp107[1], pp106[5], pp99[3], pp92[1]}, gpcOutL0_103);
gpc006 gpcL0_104 ({pp129[4], pp122[2], pp115[0], pp114[4], pp107[2], pp100[0]}, gpcOutL0_104);
gpc006 gpcL0_105 ({pp129[5], pp122[3], pp115[1], pp114[5], pp107[3], pp100[1]}, gpcOutL0_105);
gpc006 gpcL0_106 ({pp137[4], pp130[2], pp123[0], pp122[4], pp115[2], pp108[0]}, gpcOutL0_106);
gpc006 gpcL0_107 ({pp137[5], pp130[3], pp123[1], pp122[5], pp115[3], pp108[1]}, gpcOutL0_107);
gpc006 gpcL0_108 ({pp145[4], pp138[2], pp131[0], pp130[4], pp123[2], pp116[0]}, gpcOutL0_108);
gpc006 gpcL0_109 ({pp145[5], pp138[3], pp131[1], pp130[5], pp123[3], pp116[1]}, gpcOutL0_109);
gpc006 gpcL0_110 ({pp153[4], pp146[2], pp139[0], pp138[4], pp131[2], pp124[0]}, gpcOutL0_110);
gpc006 gpcL0_111 ({pp153[5], pp146[3], pp139[1], pp138[5], pp131[3], pp124[1]}, gpcOutL0_111);
gpc006 gpcL0_112 ({pp161[4], pp154[2], pp147[0], pp146[4], pp139[2], pp132[0]}, gpcOutL0_112);
gpc006 gpcL0_113 ({pp161[5], pp154[3], pp147[1], pp146[5], pp139[3], pp132[1]}, gpcOutL0_113);
gpc006 gpcL0_114 ({pp169[4], pp162[2], pp155[0], pp154[4], pp147[2], pp140[0]}, gpcOutL0_114);
gpc006 gpcL0_115 ({pp169[5], pp162[3], pp155[1], pp154[5], pp147[3], pp140[1]}, gpcOutL0_115);
gpc006 gpcL0_116 ({pp177[4], pp170[2], pp163[0], pp162[4], pp155[2], pp148[0]}, gpcOutL0_116);
gpc006 gpcL0_117 ({pp177[5], pp170[3], pp163[1], pp162[5], pp155[3], pp148[1]}, gpcOutL0_117);
gpc006 gpcL0_118 ({pp185[4], pp178[2], pp171[0], pp170[4], pp163[2], pp156[0]}, gpcOutL0_118);
gpc006 gpcL0_119 ({pp185[5], pp178[3], pp171[1], pp170[5], pp163[3], pp156[1]}, gpcOutL0_119);
gpc006 gpcL0_120 ({pp193[4], pp186[2], pp179[0], pp178[4], pp171[2], pp164[0]}, gpcOutL0_120);
gpc006 gpcL0_121 ({pp193[5], pp186[3], pp179[1], pp178[5], pp171[3], pp164[1]}, gpcOutL0_121);
gpc006 gpcL0_122 ({pp201[4], pp194[2], pp187[0], pp186[4], pp179[2], pp172[0]}, gpcOutL0_122);
gpc006 gpcL0_123 ({pp201[5], pp194[3], pp187[1], pp186[5], pp179[3], pp172[1]}, gpcOutL0_123);
gpc006 gpcL0_124 ({pp209[4], pp202[2], pp195[0], pp194[4], pp187[2], pp180[0]}, gpcOutL0_124);
gpc006 gpcL0_125 ({pp209[5], pp202[3], pp195[1], pp194[5], pp187[3], pp180[1]}, gpcOutL0_125);
gpc006 gpcL0_126 ({pp217[4], pp210[2], pp203[0], pp202[4], pp195[2], pp188[0]}, gpcOutL0_126);
gpc006 gpcL0_127 ({pp217[5], pp210[3], pp203[1], pp202[5], pp195[3], pp188[1]}, gpcOutL0_127);
gpc006 gpcL0_128 ({pp218[2], pp211[0], pp210[4], pp203[2], pp196[0], pp195[4]}, gpcOutL0_128);
gpc006 gpcL0_129 ({pp218[3], pp211[1], pp210[5], pp203[3], pp196[1], pp195[5]}, gpcOutL0_129);
gpc006 gpcL0_130 ({pp219[0], pp218[4], pp211[2], pp204[0], pp203[4], pp196[2]}, gpcOutL0_130);
gpc006 gpcL0_131 ({pp219[1], pp218[5], pp211[3], pp204[1], pp203[5], pp196[3]}, gpcOutL0_131);
gpc006 gpcL0_132 ({pp219[2], pp212[0], pp211[4], pp204[2], pp197[0], pp196[4]}, gpcOutL0_132);
gpc006 gpcL0_133 ({pp219[3], pp212[1], pp211[5], pp204[3], pp197[1], pp196[5]}, gpcOutL0_133);
gpc006 gpcL0_134 ({pp220[0], pp219[4], pp212[2], pp205[0], pp204[4], pp197[2]}, gpcOutL0_134);
gpc006 gpcL0_135 ({pp220[1], pp219[5], pp212[3], pp205[1], pp204[5], pp197[3]}, gpcOutL0_135);
gpc006 gpcL0_136 ({pp220[2], pp213[0], pp212[4], pp205[2], pp198[0], pp197[4]}, gpcOutL0_136);
gpc006 gpcL0_137 ({pp220[3], pp213[1], pp212[5], pp205[3], pp198[1], pp197[5]}, gpcOutL0_137);
gpc006 gpcL0_138 ({pp221[0], pp220[4], pp213[2], pp206[0], pp205[4], pp198[2]}, gpcOutL0_138);
gpc006 gpcL0_139 ({pp221[1], pp220[5], pp213[3], pp206[1], pp205[5], pp198[3]}, gpcOutL0_139);
gpc006 gpcL0_140 ({pp221[2], pp214[0], pp213[4], pp206[2], pp199[0], pp198[4]}, gpcOutL0_140);
gpc006 gpcL0_141 ({pp221[3], pp214[1], pp213[5], pp206[3], pp199[1], pp198[5]}, gpcOutL0_141);
gpc006 gpcL0_142 ({pp222[0], pp221[4], pp214[2], pp207[0], pp206[4], pp199[2]}, gpcOutL0_142);
gpc006 gpcL0_143 ({pp222[1], pp221[5], pp214[3], pp207[1], pp206[5], pp199[3]}, gpcOutL0_143);
gpc006 gpcL0_144 ({pp35[4], pp28[2], pp21[0], pp20[4], pp13[2], pp6[0]}, gpcOutL0_144);
gpc006 gpcL0_145 ({pp35[5], pp28[3], pp21[1], pp20[5], pp13[3], pp6[1]}, gpcOutL0_145);
gpc006 gpcL0_146 ({pp43[4], pp36[2], pp29[0], pp28[4], pp21[2], pp14[0]}, gpcOutL0_146);
gpc006 gpcL0_147 ({pp43[5], pp36[3], pp29[1], pp28[5], pp21[3], pp14[1]}, gpcOutL0_147);
gpc006 gpcL0_148 ({pp51[4], pp44[2], pp37[0], pp36[4], pp29[2], pp22[0]}, gpcOutL0_148);
gpc006 gpcL0_149 ({pp51[5], pp44[3], pp37[1], pp36[5], pp29[3], pp22[1]}, gpcOutL0_149);
gpc006 gpcL0_150 ({pp59[4], pp52[2], pp45[0], pp44[4], pp37[2], pp30[0]}, gpcOutL0_150);
gpc006 gpcL0_151 ({pp59[5], pp52[3], pp45[1], pp44[5], pp37[3], pp30[1]}, gpcOutL0_151);
gpc006 gpcL0_152 ({pp67[4], pp60[2], pp53[0], pp52[4], pp45[2], pp38[0]}, gpcOutL0_152);
gpc006 gpcL0_153 ({pp67[5], pp60[3], pp53[1], pp52[5], pp45[3], pp38[1]}, gpcOutL0_153);
gpc006 gpcL0_154 ({pp75[4], pp68[2], pp61[0], pp60[4], pp53[2], pp46[0]}, gpcOutL0_154);
gpc006 gpcL0_155 ({pp75[5], pp68[3], pp61[1], pp60[5], pp53[3], pp46[1]}, gpcOutL0_155);
gpc006 gpcL0_156 ({pp83[4], pp76[2], pp69[0], pp68[4], pp61[2], pp54[0]}, gpcOutL0_156);
gpc006 gpcL0_157 ({pp83[5], pp76[3], pp69[1], pp68[5], pp61[3], pp54[1]}, gpcOutL0_157);
gpc006 gpcL0_158 ({pp91[4], pp84[2], pp77[0], pp76[4], pp69[2], pp62[0]}, gpcOutL0_158);
gpc006 gpcL0_159 ({pp91[5], pp84[3], pp77[1], pp76[5], pp69[3], pp62[1]}, gpcOutL0_159);
gpc006 gpcL0_160 ({pp99[4], pp92[2], pp85[0], pp84[4], pp77[2], pp70[0]}, gpcOutL0_160);
gpc006 gpcL0_161 ({pp99[5], pp92[3], pp85[1], pp84[5], pp77[3], pp70[1]}, gpcOutL0_161);
gpc006 gpcL0_162 ({pp107[4], pp100[2], pp93[0], pp92[4], pp85[2], pp78[0]}, gpcOutL0_162);
gpc006 gpcL0_163 ({pp107[5], pp100[3], pp93[1], pp92[5], pp85[3], pp78[1]}, gpcOutL0_163);
gpc006 gpcL0_164 ({pp115[4], pp108[2], pp101[0], pp100[4], pp93[2], pp86[0]}, gpcOutL0_164);
gpc006 gpcL0_165 ({pp115[5], pp108[3], pp101[1], pp100[5], pp93[3], pp86[1]}, gpcOutL0_165);
gpc006 gpcL0_166 ({pp123[4], pp116[2], pp109[0], pp108[4], pp101[2], pp94[0]}, gpcOutL0_166);
gpc006 gpcL0_167 ({pp123[5], pp116[3], pp109[1], pp108[5], pp101[3], pp94[1]}, gpcOutL0_167);
gpc006 gpcL0_168 ({pp131[4], pp124[2], pp117[0], pp116[4], pp109[2], pp102[0]}, gpcOutL0_168);
gpc006 gpcL0_169 ({pp131[5], pp124[3], pp117[1], pp116[5], pp109[3], pp102[1]}, gpcOutL0_169);
gpc006 gpcL0_170 ({pp139[4], pp132[2], pp125[0], pp124[4], pp117[2], pp110[0]}, gpcOutL0_170);
gpc006 gpcL0_171 ({pp139[5], pp132[3], pp125[1], pp124[5], pp117[3], pp110[1]}, gpcOutL0_171);
gpc006 gpcL0_172 ({pp147[4], pp140[2], pp133[0], pp132[4], pp125[2], pp118[0]}, gpcOutL0_172);
gpc006 gpcL0_173 ({pp147[5], pp140[3], pp133[1], pp132[5], pp125[3], pp118[1]}, gpcOutL0_173);
gpc006 gpcL0_174 ({pp155[4], pp148[2], pp141[0], pp140[4], pp133[2], pp126[0]}, gpcOutL0_174);
gpc006 gpcL0_175 ({pp155[5], pp148[3], pp141[1], pp140[5], pp133[3], pp126[1]}, gpcOutL0_175);
gpc006 gpcL0_176 ({pp163[4], pp156[2], pp149[0], pp148[4], pp141[2], pp134[0]}, gpcOutL0_176);
gpc006 gpcL0_177 ({pp163[5], pp156[3], pp149[1], pp148[5], pp141[3], pp134[1]}, gpcOutL0_177);
gpc006 gpcL0_178 ({pp171[4], pp164[2], pp157[0], pp156[4], pp149[2], pp142[0]}, gpcOutL0_178);
gpc006 gpcL0_179 ({pp171[5], pp164[3], pp157[1], pp156[5], pp149[3], pp142[1]}, gpcOutL0_179);
gpc006 gpcL0_180 ({pp179[4], pp172[2], pp165[0], pp164[4], pp157[2], pp150[0]}, gpcOutL0_180);
gpc006 gpcL0_181 ({pp179[5], pp172[3], pp165[1], pp164[5], pp157[3], pp150[1]}, gpcOutL0_181);
gpc006 gpcL0_182 ({pp187[4], pp180[2], pp173[0], pp172[4], pp165[2], pp158[0]}, gpcOutL0_182);
gpc006 gpcL0_183 ({pp187[5], pp180[3], pp173[1], pp172[5], pp165[3], pp158[1]}, gpcOutL0_183);
gpc006 gpcL0_184 ({pp188[2], pp181[0], pp180[4], pp173[2], pp166[0], pp165[4]}, gpcOutL0_184);
gpc006 gpcL0_185 ({pp188[3], pp181[1], pp180[5], pp173[3], pp166[1], pp165[5]}, gpcOutL0_185);
gpc006 gpcL0_186 ({pp189[0], pp188[4], pp181[2], pp174[0], pp173[4], pp166[2]}, gpcOutL0_186);
gpc006 gpcL0_187 ({pp189[1], pp188[5], pp181[3], pp174[1], pp173[5], pp166[3]}, gpcOutL0_187);
gpc006 gpcL0_188 ({pp189[2], pp182[0], pp181[4], pp174[2], pp167[0], pp166[4]}, gpcOutL0_188);
gpc006 gpcL0_189 ({pp189[3], pp182[1], pp181[5], pp174[3], pp167[1], pp166[5]}, gpcOutL0_189);
gpc006 gpcL0_190 ({pp190[0], pp189[4], pp182[2], pp175[0], pp174[4], pp167[2]}, gpcOutL0_190);
gpc006 gpcL0_191 ({pp190[1], pp189[5], pp182[3], pp175[1], pp174[5], pp167[3]}, gpcOutL0_191);
gpc006 gpcL0_192 ({pp37[4], pp30[2], pp23[0], pp22[4], pp15[2], pp7[4]}, gpcOutL0_192);
gpc006 gpcL0_193 ({pp37[5], pp30[3], pp23[1], pp22[5], pp15[3], pp7[5]}, gpcOutL0_193);
gpc006 gpcL0_194 ({pp45[4], pp38[2], pp31[0], pp30[4], pp23[2], pp15[4]}, gpcOutL0_194);
gpc006 gpcL0_195 ({pp45[5], pp38[3], pp31[1], pp30[5], pp23[3], pp15[5]}, gpcOutL0_195);
gpc006 gpcL0_196 ({pp53[4], pp46[2], pp39[0], pp38[4], pp31[2], pp23[4]}, gpcOutL0_196);
gpc006 gpcL0_197 ({pp53[5], pp46[3], pp39[1], pp38[5], pp31[3], pp23[5]}, gpcOutL0_197);
gpc006 gpcL0_198 ({pp61[4], pp54[2], pp47[0], pp46[4], pp39[2], pp31[4]}, gpcOutL0_198);
gpc006 gpcL0_199 ({pp61[5], pp54[3], pp47[1], pp46[5], pp39[3], pp31[5]}, gpcOutL0_199);
gpc006 gpcL0_200 ({pp69[4], pp62[2], pp55[0], pp54[4], pp47[2], pp39[4]}, gpcOutL0_200);
gpc006 gpcL0_201 ({pp69[5], pp62[3], pp55[1], pp54[5], pp47[3], pp39[5]}, gpcOutL0_201);
gpc006 gpcL0_202 ({pp77[4], pp70[2], pp63[0], pp62[4], pp55[2], pp47[4]}, gpcOutL0_202);
gpc006 gpcL0_203 ({pp77[5], pp70[3], pp63[1], pp62[5], pp55[3], pp47[5]}, gpcOutL0_203);
gpc006 gpcL0_204 ({pp85[4], pp78[2], pp71[0], pp70[4], pp63[2], pp55[4]}, gpcOutL0_204);
gpc006 gpcL0_205 ({pp85[5], pp78[3], pp71[1], pp70[5], pp63[3], pp55[5]}, gpcOutL0_205);
gpc006 gpcL0_206 ({pp93[4], pp86[2], pp79[0], pp78[4], pp71[2], pp63[4]}, gpcOutL0_206);
gpc006 gpcL0_207 ({pp93[5], pp86[3], pp79[1], pp78[5], pp71[3], pp63[5]}, gpcOutL0_207);
gpc006 gpcL0_208 ({pp101[4], pp94[2], pp87[0], pp86[4], pp79[2], pp71[4]}, gpcOutL0_208);
gpc006 gpcL0_209 ({pp101[5], pp94[3], pp87[1], pp86[5], pp79[3], pp71[5]}, gpcOutL0_209);
gpc006 gpcL0_210 ({pp109[4], pp102[2], pp95[0], pp94[4], pp87[2], pp79[4]}, gpcOutL0_210);
gpc006 gpcL0_211 ({pp109[5], pp102[3], pp95[1], pp94[5], pp87[3], pp79[5]}, gpcOutL0_211);
gpc006 gpcL0_212 ({pp117[4], pp110[2], pp103[0], pp102[4], pp95[2], pp87[4]}, gpcOutL0_212);
gpc006 gpcL0_213 ({pp117[5], pp110[3], pp103[1], pp102[5], pp95[3], pp87[5]}, gpcOutL0_213);
gpc006 gpcL0_214 ({pp125[4], pp118[2], pp111[0], pp110[4], pp103[2], pp95[4]}, gpcOutL0_214);
gpc006 gpcL0_215 ({pp125[5], pp118[3], pp111[1], pp110[5], pp103[3], pp95[5]}, gpcOutL0_215);
gpc006 gpcL0_216 ({pp133[4], pp126[2], pp119[0], pp118[4], pp111[2], pp103[4]}, gpcOutL0_216);
gpc006 gpcL0_217 ({pp133[5], pp126[3], pp119[1], pp118[5], pp111[3], pp103[5]}, gpcOutL0_217);
gpc006 gpcL0_218 ({pp141[4], pp134[2], pp127[0], pp126[4], pp119[2], pp111[4]}, gpcOutL0_218);
gpc006 gpcL0_219 ({pp141[5], pp134[3], pp127[1], pp126[5], pp119[3], pp111[5]}, gpcOutL0_219);
gpc006 gpcL0_220 ({pp149[4], pp142[2], pp135[0], pp134[4], pp127[2], pp119[4]}, gpcOutL0_220);
gpc006 gpcL0_221 ({pp149[5], pp142[3], pp135[1], pp134[5], pp127[3], pp119[5]}, gpcOutL0_221);
gpc006 gpcL0_222 ({pp157[4], pp150[2], pp143[0], pp142[4], pp135[2], pp127[4]}, gpcOutL0_222);
gpc006 gpcL0_223 ({pp157[5], pp150[3], pp143[1], pp142[5], pp135[3], pp127[5]}, gpcOutL0_223);
gpc015 gpcL0_224 ({pp24[1], pp24[0], pp16[2], pp9[0], pp8[4], pp1[2]}, gpcOutL0_224);
gpc015 gpcL0_225 ({pp25[5], pp25[4], pp18[2], pp11[0], pp10[4], pp3[2]}, gpcOutL0_225);
gpc015 gpcL0_226 ({pp27[5], pp27[4], pp20[2], pp13[0], pp12[4], pp5[2]}, gpcOutL0_226);
gpc015 gpcL0_227 ({pp29[5], pp29[4], pp22[2], pp15[0], pp14[4], pp7[2]}, gpcOutL0_227);
gpc015 gpcL0_228 ({pp158[3], pp158[2], pp151[0], pp150[4], pp143[2], pp135[4]}, gpcOutL0_228);
gpc015 gpcL0_229 ({pp190[3], pp190[2], pp183[0], pp182[4], pp175[2], pp167[4]}, gpcOutL0_229);
gpc015 gpcL0_230 ({pp222[3], pp222[2], pp215[0], pp214[4], pp207[2], pp199[4]}, gpcOutL0_230);
gpc015 gpcL0_231 ({pp254[3], pp254[2], pp247[0], pp246[4], pp239[2], pp231[4]}, gpcOutL0_231);
gpc014 gpcL0_232 ({pp16[1], pp16[0], pp8[2], pp1[0], pp0[4]}, gpcOutL0_232);
gpc014 gpcL0_233 ({pp1[4], pp16[3], pp9[1], pp8[5], pp1[3]}, gpcOutL0_233);
gpc014 gpcL0_234 ({pp17[5], pp17[4], pp10[2], pp3[0], pp2[4]}, gpcOutL0_234);
gpc014 gpcL0_235 ({pp3[4], pp18[3], pp11[1], pp10[5], pp3[3]}, gpcOutL0_235);
gpc014 gpcL0_236 ({pp19[5], pp19[4], pp12[2], pp5[0], pp4[4]}, gpcOutL0_236);
gpc014 gpcL0_237 ({pp5[4], pp20[3], pp13[1], pp12[5], pp5[3]}, gpcOutL0_237);
gpc014 gpcL0_238 ({pp21[5], pp21[4], pp14[2], pp7[0], pp6[4]}, gpcOutL0_238);
gpc014 gpcL0_239 ({pp159[0], pp151[1], pp150[5], pp143[3], pp135[5]}, gpcOutL0_239);
gpc014 gpcL0_240 ({pp159[2], pp159[1], pp158[5], pp151[3], pp143[5]}, gpcOutL0_240);
gpc014 gpcL0_241 ({pp191[0], pp183[1], pp182[5], pp175[3], pp167[5]}, gpcOutL0_241);
gpc014 gpcL0_242 ({pp191[2], pp191[1], pp190[5], pp183[3], pp175[5]}, gpcOutL0_242);
gpc014 gpcL0_243 ({pp223[0], pp215[1], pp214[5], pp207[3], pp199[5]}, gpcOutL0_243);
gpc014 gpcL0_244 ({pp223[2], pp223[1], pp222[5], pp215[3], pp207[5]}, gpcOutL0_244);
gpc014 gpcL0_245 ({pp255[0], pp247[1], pp246[5], pp239[3], pp231[5]}, gpcOutL0_245);
gpc014 gpcL0_246 ({pp255[2], pp255[1], pp254[5], pp247[3], pp239[5]}, gpcOutL0_246);
gpc003 gpcL0_247 ({pp8[3], pp1[1], pp0[5]}, gpcOutL0_247);
gpc003 gpcL0_248 ({pp10[3], pp3[1], pp2[5]}, gpcOutL0_248);
gpc003 gpcL0_249 ({pp12[3], pp5[1], pp4[5]}, gpcOutL0_249);
gpc003 gpcL0_250 ({pp14[3], pp7[1], pp6[5]}, gpcOutL0_250);
gpc003 gpcL0_251 ({pp22[3], pp15[1], pp14[5]}, gpcOutL0_251);
gpc003 gpcL0_252 ({pp158[4], pp151[2], pp143[4]}, gpcOutL0_252);
gpc003 gpcL0_253 ({pp190[4], pp183[2], pp175[4]}, gpcOutL0_253);
gpc003 gpcL0_254 ({pp222[4], pp215[2], pp207[4]}, gpcOutL0_254);
gpc003 gpcL0_255 ({pp254[4], pp247[2], pp239[4]}, gpcOutL0_255);
gpc022 gpcL0_256 ({pp9[5], pp2[3], pp9[4], pp2[2]}, gpcOutL0_256);
gpc022 gpcL0_257 ({pp11[5], pp4[3], pp11[4], pp4[2]}, gpcOutL0_257);
gpc022 gpcL0_258 ({pp13[5], pp6[3], pp13[4], pp6[2]}, gpcOutL0_258);
gpc022 gpcL0_259 ({pp8[1], pp0[3], pp8[0], pp0[2]}, gpcOutL0_259);

// level 1
wire [2:0]  gpcOutL1_0;
wire [2:0]  gpcOutL1_1;
wire [2:0]  gpcOutL1_2;
wire [2:0]  gpcOutL1_3;
wire [2:0]  gpcOutL1_4;
wire [2:0]  gpcOutL1_5;
wire [2:0]  gpcOutL1_6;
wire [2:0]  gpcOutL1_7;
wire [2:0]  gpcOutL1_8;
wire [2:0]  gpcOutL1_9;
wire [2:0]  gpcOutL1_10;
wire [2:0]  gpcOutL1_11;
wire [2:0]  gpcOutL1_12;
wire [2:0]  gpcOutL1_13;
wire [2:0]  gpcOutL1_14;
wire [2:0]  gpcOutL1_15;
wire [2:0]  gpcOutL1_16;
wire [2:0]  gpcOutL1_17;
wire [2:0]  gpcOutL1_18;
wire [2:0]  gpcOutL1_19;
wire [2:0]  gpcOutL1_20;
wire [2:0]  gpcOutL1_21;
wire [2:0]  gpcOutL1_22;
wire [2:0]  gpcOutL1_23;
wire [2:0]  gpcOutL1_24;
wire [2:0]  gpcOutL1_25;
wire [2:0]  gpcOutL1_26;
wire [2:0]  gpcOutL1_27;
wire [2:0]  gpcOutL1_28;
wire [2:0]  gpcOutL1_29;
wire [2:0]  gpcOutL1_30;
wire [2:0]  gpcOutL1_31;
wire [2:0]  gpcOutL1_32;
wire [2:0]  gpcOutL1_33;
wire [2:0]  gpcOutL1_34;
wire [2:0]  gpcOutL1_35;
wire [2:0]  gpcOutL1_36;
wire [2:0]  gpcOutL1_37;
wire [2:0]  gpcOutL1_38;
wire [2:0]  gpcOutL1_39;
wire [2:0]  gpcOutL1_40;
wire [2:0]  gpcOutL1_41;
wire [2:0]  gpcOutL1_42;
wire [2:0]  gpcOutL1_43;
wire [2:0]  gpcOutL1_44;
wire [2:0]  gpcOutL1_45;
wire [2:0]  gpcOutL1_46;
wire [2:0]  gpcOutL1_47;
wire [2:0]  gpcOutL1_48;
wire [2:0]  gpcOutL1_49;
wire [2:0]  gpcOutL1_50;
wire [2:0]  gpcOutL1_51;
wire [2:0]  gpcOutL1_52;
wire [2:0]  gpcOutL1_53;
wire [2:0]  gpcOutL1_54;
wire [2:0]  gpcOutL1_55;
wire [2:0]  gpcOutL1_56;
wire [2:0]  gpcOutL1_57;
wire [2:0]  gpcOutL1_58;
wire [2:0]  gpcOutL1_59;
wire [2:0]  gpcOutL1_60;
wire [2:0]  gpcOutL1_61;
wire [2:0]  gpcOutL1_62;
wire [2:0]  gpcOutL1_63;
wire [2:0]  gpcOutL1_64;
wire [2:0]  gpcOutL1_65;
wire [2:0]  gpcOutL1_66;
wire [2:0]  gpcOutL1_67;
wire [2:0]  gpcOutL1_68;
wire [2:0]  gpcOutL1_69;
wire [2:0]  gpcOutL1_70;
wire [2:0]  gpcOutL1_71;
wire [2:0]  gpcOutL1_72;
wire [2:0]  gpcOutL1_73;
wire [2:0]  gpcOutL1_74;
wire [2:0]  gpcOutL1_75;
wire [2:0]  gpcOutL1_76;
wire [2:0]  gpcOutL1_77;
wire [2:0]  gpcOutL1_78;
wire [2:0]  gpcOutL1_79;
wire [2:0]  gpcOutL1_80;
wire [2:0]  gpcOutL1_81;
wire [2:0]  gpcOutL1_82;
wire [2:0]  gpcOutL1_83;
wire [2:0]  gpcOutL1_84;
wire [2:0]  gpcOutL1_85;
wire [2:0]  gpcOutL1_86;
wire [2:0]  gpcOutL1_87;
wire [2:0]  gpcOutL1_88;
wire [2:0]  gpcOutL1_89;
wire [2:0]  gpcOutL1_90;
wire [2:0]  gpcOutL1_91;
wire [2:0]  gpcOutL1_92;
wire [2:0]  gpcOutL1_93;
wire [2:0]  gpcOutL1_94;
wire [2:0]  gpcOutL1_95;
wire [2:0]  gpcOutL1_96;
wire [2:0]  gpcOutL1_97;
wire [2:0]  gpcOutL1_98;
wire [2:0]  gpcOutL1_99;
wire [2:0]  gpcOutL1_100;
wire [2:0]  gpcOutL1_101;
wire [2:0]  gpcOutL1_102;
wire [2:0]  gpcOutL1_103;
wire [2:0]  gpcOutL1_104;
wire [2:0]  gpcOutL1_105;
wire [2:0]  gpcOutL1_106;
wire [2:0]  gpcOutL1_107;
wire [2:0]  gpcOutL1_108;
wire [2:0]  gpcOutL1_109;
wire [2:0]  gpcOutL1_110;
wire [2:0]  gpcOutL1_111;
wire [2:0]  gpcOutL1_112;
wire [2:0]  gpcOutL1_113;
wire [2:0]  gpcOutL1_114;
wire [2:0]  gpcOutL1_115;
wire [2:0]  gpcOutL1_116;
wire [2:0]  gpcOutL1_117;
wire [2:0]  gpcOutL1_118;
wire [2:0]  gpcOutL1_119;
wire [2:0]  gpcOutL1_120;
wire [2:0]  gpcOutL1_121;
wire [2:0]  gpcOutL1_122;
wire [2:0]  gpcOutL1_123;
wire [2:0]  gpcOutL1_124;
wire [2:0]  gpcOutL1_125;
wire [2:0]  gpcOutL1_126;
wire [1:0]  gpcOutL1_127;
wire [1:0]  gpcOutL1_128;
wire [1:0]  gpcOutL1_129;
wire [1:0]  gpcOutL1_130;
wire [1:0]  gpcOutL1_131;
wire [2:0]  gpcOutL1_132;
wire [3:0]  gpcOutL1_133;

gpc006 gpcL1_0 ({gpcOutL0_248[1], gpcOutL0_234[2], gpcOutL0_225[0], gpcOutL0_6[0], gpcOutL0_5[1], gpcOutL0_4[2]}, gpcOutL1_0);
gpc006 gpcL1_1 ({gpcOutL0_235[1], gpcOutL0_225[2], gpcOutL0_80[0], gpcOutL0_8[0], gpcOutL0_7[1], gpcOutL0_6[2]}, gpcOutL1_1);
gpc006 gpcL1_2 ({gpcOutL0_235[2], gpcOutL0_81[0], gpcOutL0_80[1], gpcOutL0_9[0], gpcOutL0_8[1], gpcOutL0_7[2]}, gpcOutL1_2);
gpc006 gpcL1_3 ({gpcOutL0_257[0], gpcOutL0_82[0], gpcOutL0_81[1], gpcOutL0_80[2], gpcOutL0_10[0], gpcOutL0_9[1]}, gpcOutL1_3);
gpc006 gpcL1_4 ({gpcOutL0_257[1], gpcOutL0_83[0], gpcOutL0_82[1], gpcOutL0_81[2], gpcOutL0_11[0], gpcOutL0_10[1]}, gpcOutL1_4);
gpc006 gpcL1_5 ({gpcOutL0_257[2], gpcOutL0_236[0], gpcOutL0_84[0], gpcOutL0_83[1], gpcOutL0_82[2], gpcOutL0_12[0]}, gpcOutL1_5);
gpc006 gpcL1_6 ({gpcOutL0_249[0], gpcOutL0_236[1], gpcOutL0_85[0], gpcOutL0_84[1], gpcOutL0_83[2], gpcOutL0_13[0]}, gpcOutL1_6);
gpc006 gpcL1_7 ({gpcOutL0_249[1], gpcOutL0_236[2], gpcOutL0_226[0], gpcOutL0_86[0], gpcOutL0_85[1], gpcOutL0_84[2]}, gpcOutL1_7);
gpc006 gpcL1_8 ({gpcOutL0_237[0], gpcOutL0_226[1], gpcOutL0_87[0], gpcOutL0_86[1], gpcOutL0_85[2], gpcOutL0_15[0]}, gpcOutL1_8);
gpc006 gpcL1_9 ({gpcOutL0_237[1], gpcOutL0_226[2], gpcOutL0_144[0], gpcOutL0_88[0], gpcOutL0_87[1], gpcOutL0_86[2]}, gpcOutL1_9);
gpc006 gpcL1_10 ({gpcOutL0_237[2], gpcOutL0_145[0], gpcOutL0_144[1], gpcOutL0_89[0], gpcOutL0_88[1], gpcOutL0_87[2]}, gpcOutL1_10);
gpc006 gpcL1_11 ({gpcOutL0_258[0], gpcOutL0_146[0], gpcOutL0_145[1], gpcOutL0_144[2], gpcOutL0_90[0], gpcOutL0_89[1]}, gpcOutL1_11);
gpc006 gpcL1_12 ({gpcOutL0_258[1], gpcOutL0_147[0], gpcOutL0_146[1], gpcOutL0_145[2], gpcOutL0_91[0], gpcOutL0_90[1]}, gpcOutL1_12);
gpc006 gpcL1_13 ({gpcOutL0_258[2], gpcOutL0_238[0], gpcOutL0_148[0], gpcOutL0_147[1], gpcOutL0_146[2], gpcOutL0_92[0]}, gpcOutL1_13);
gpc006 gpcL1_14 ({gpcOutL0_250[0], gpcOutL0_238[1], gpcOutL0_149[0], gpcOutL0_148[1], gpcOutL0_147[2], gpcOutL0_93[0]}, gpcOutL1_14);
gpc006 gpcL1_15 ({gpcOutL0_250[1], gpcOutL0_238[2], gpcOutL0_227[0], gpcOutL0_150[0], gpcOutL0_149[1], gpcOutL0_148[2]}, gpcOutL1_15);
gpc006 gpcL1_16 ({gpcOutL0_251[0], gpcOutL0_227[1], gpcOutL0_151[0], gpcOutL0_150[1], gpcOutL0_149[2], gpcOutL0_95[0]}, gpcOutL1_16);
gpc006 gpcL1_17 ({gpcOutL0_251[1], gpcOutL0_227[2], gpcOutL0_192[0], gpcOutL0_152[0], gpcOutL0_151[1], gpcOutL0_150[2]}, gpcOutL1_17);
gpc006 gpcL1_18 ({gpcOutL0_193[0], gpcOutL0_192[1], gpcOutL0_153[0], gpcOutL0_152[1], gpcOutL0_151[2], gpcOutL0_97[0]}, gpcOutL1_18);
gpc006 gpcL1_19 ({gpcOutL0_194[0], gpcOutL0_193[1], gpcOutL0_192[2], gpcOutL0_154[0], gpcOutL0_153[1], gpcOutL0_152[2]}, gpcOutL1_19);
gpc006 gpcL1_20 ({gpcOutL0_195[0], gpcOutL0_194[1], gpcOutL0_193[2], gpcOutL0_155[0], gpcOutL0_154[1], gpcOutL0_153[2]}, gpcOutL1_20);
gpc006 gpcL1_21 ({gpcOutL0_196[0], gpcOutL0_195[1], gpcOutL0_194[2], gpcOutL0_156[0], gpcOutL0_155[1], gpcOutL0_154[2]}, gpcOutL1_21);
gpc006 gpcL1_22 ({gpcOutL0_197[0], gpcOutL0_196[1], gpcOutL0_195[2], gpcOutL0_157[0], gpcOutL0_156[1], gpcOutL0_155[2]}, gpcOutL1_22);
gpc006 gpcL1_23 ({gpcOutL0_198[0], gpcOutL0_197[1], gpcOutL0_196[2], gpcOutL0_158[0], gpcOutL0_157[1], gpcOutL0_156[2]}, gpcOutL1_23);
gpc006 gpcL1_24 ({gpcOutL0_199[0], gpcOutL0_198[1], gpcOutL0_197[2], gpcOutL0_159[0], gpcOutL0_158[1], gpcOutL0_157[2]}, gpcOutL1_24);
gpc006 gpcL1_25 ({gpcOutL0_200[0], gpcOutL0_199[1], gpcOutL0_198[2], gpcOutL0_160[0], gpcOutL0_159[1], gpcOutL0_158[2]}, gpcOutL1_25);
gpc006 gpcL1_26 ({gpcOutL0_201[0], gpcOutL0_200[1], gpcOutL0_199[2], gpcOutL0_161[0], gpcOutL0_160[1], gpcOutL0_159[2]}, gpcOutL1_26);
gpc006 gpcL1_27 ({gpcOutL0_202[0], gpcOutL0_201[1], gpcOutL0_200[2], gpcOutL0_162[0], gpcOutL0_161[1], gpcOutL0_160[2]}, gpcOutL1_27);
gpc006 gpcL1_28 ({gpcOutL0_203[0], gpcOutL0_202[1], gpcOutL0_201[2], gpcOutL0_163[0], gpcOutL0_162[1], gpcOutL0_161[2]}, gpcOutL1_28);
gpc006 gpcL1_29 ({gpcOutL0_204[0], gpcOutL0_203[1], gpcOutL0_202[2], gpcOutL0_164[0], gpcOutL0_163[1], gpcOutL0_162[2]}, gpcOutL1_29);
gpc006 gpcL1_30 ({gpcOutL0_205[0], gpcOutL0_204[1], gpcOutL0_203[2], gpcOutL0_165[0], gpcOutL0_164[1], gpcOutL0_163[2]}, gpcOutL1_30);
gpc006 gpcL1_31 ({gpcOutL0_206[0], gpcOutL0_205[1], gpcOutL0_204[2], gpcOutL0_166[0], gpcOutL0_165[1], gpcOutL0_164[2]}, gpcOutL1_31);
gpc006 gpcL1_32 ({gpcOutL0_207[0], gpcOutL0_206[1], gpcOutL0_205[2], gpcOutL0_167[0], gpcOutL0_166[1], gpcOutL0_165[2]}, gpcOutL1_32);
gpc006 gpcL1_33 ({gpcOutL0_208[0], gpcOutL0_207[1], gpcOutL0_206[2], gpcOutL0_168[0], gpcOutL0_167[1], gpcOutL0_166[2]}, gpcOutL1_33);
gpc006 gpcL1_34 ({gpcOutL0_209[0], gpcOutL0_208[1], gpcOutL0_207[2], gpcOutL0_169[0], gpcOutL0_168[1], gpcOutL0_167[2]}, gpcOutL1_34);
gpc006 gpcL1_35 ({gpcOutL0_210[0], gpcOutL0_209[1], gpcOutL0_208[2], gpcOutL0_170[0], gpcOutL0_169[1], gpcOutL0_168[2]}, gpcOutL1_35);
gpc006 gpcL1_36 ({gpcOutL0_211[0], gpcOutL0_210[1], gpcOutL0_209[2], gpcOutL0_171[0], gpcOutL0_170[1], gpcOutL0_169[2]}, gpcOutL1_36);
gpc006 gpcL1_37 ({gpcOutL0_212[0], gpcOutL0_211[1], gpcOutL0_210[2], gpcOutL0_172[0], gpcOutL0_171[1], gpcOutL0_170[2]}, gpcOutL1_37);
gpc006 gpcL1_38 ({gpcOutL0_213[0], gpcOutL0_212[1], gpcOutL0_211[2], gpcOutL0_173[0], gpcOutL0_172[1], gpcOutL0_171[2]}, gpcOutL1_38);
gpc006 gpcL1_39 ({gpcOutL0_214[0], gpcOutL0_213[1], gpcOutL0_212[2], gpcOutL0_174[0], gpcOutL0_173[1], gpcOutL0_172[2]}, gpcOutL1_39);
gpc006 gpcL1_40 ({gpcOutL0_215[0], gpcOutL0_214[1], gpcOutL0_213[2], gpcOutL0_175[0], gpcOutL0_174[1], gpcOutL0_173[2]}, gpcOutL1_40);
gpc006 gpcL1_41 ({gpcOutL0_216[0], gpcOutL0_215[1], gpcOutL0_214[2], gpcOutL0_176[0], gpcOutL0_175[1], gpcOutL0_174[2]}, gpcOutL1_41);
gpc006 gpcL1_42 ({gpcOutL0_217[0], gpcOutL0_216[1], gpcOutL0_215[2], gpcOutL0_177[0], gpcOutL0_176[1], gpcOutL0_175[2]}, gpcOutL1_42);
gpc006 gpcL1_43 ({gpcOutL0_218[0], gpcOutL0_217[1], gpcOutL0_216[2], gpcOutL0_178[0], gpcOutL0_177[1], gpcOutL0_176[2]}, gpcOutL1_43);
gpc006 gpcL1_44 ({gpcOutL0_219[0], gpcOutL0_218[1], gpcOutL0_217[2], gpcOutL0_179[0], gpcOutL0_178[1], gpcOutL0_177[2]}, gpcOutL1_44);
gpc006 gpcL1_45 ({gpcOutL0_220[0], gpcOutL0_219[1], gpcOutL0_218[2], gpcOutL0_180[0], gpcOutL0_179[1], gpcOutL0_178[2]}, gpcOutL1_45);
gpc006 gpcL1_46 ({gpcOutL0_221[0], gpcOutL0_220[1], gpcOutL0_219[2], gpcOutL0_181[0], gpcOutL0_180[1], gpcOutL0_179[2]}, gpcOutL1_46);
gpc006 gpcL1_47 ({gpcOutL0_222[0], gpcOutL0_221[1], gpcOutL0_220[2], gpcOutL0_182[0], gpcOutL0_181[1], gpcOutL0_180[2]}, gpcOutL1_47);
gpc006 gpcL1_48 ({gpcOutL0_223[0], gpcOutL0_222[1], gpcOutL0_221[2], gpcOutL0_183[0], gpcOutL0_182[1], gpcOutL0_181[2]}, gpcOutL1_48);
gpc006 gpcL1_49 ({gpcOutL0_228[0], gpcOutL0_223[1], gpcOutL0_222[2], gpcOutL0_184[0], gpcOutL0_183[1], gpcOutL0_182[2]}, gpcOutL1_49);
gpc006 gpcL1_50 ({gpcOutL0_239[0], gpcOutL0_228[1], gpcOutL0_223[2], gpcOutL0_185[0], gpcOutL0_184[1], gpcOutL0_183[2]}, gpcOutL1_50);
gpc006 gpcL1_51 ({gpcOutL0_252[0], gpcOutL0_239[1], gpcOutL0_228[2], gpcOutL0_186[0], gpcOutL0_185[1], gpcOutL0_184[2]}, gpcOutL1_51);
gpc006 gpcL1_52 ({gpcOutL0_252[1], gpcOutL0_240[0], gpcOutL0_239[2], gpcOutL0_187[0], gpcOutL0_186[1], gpcOutL0_185[2]}, gpcOutL1_52);
gpc006 gpcL1_53 ({gpcOutL0_240[1], gpcOutL0_188[0], gpcOutL0_187[1], gpcOutL0_186[2], gpcOutL0_132[0], gpcOutL0_131[1]}, gpcOutL1_53);
gpc006 gpcL1_54 ({gpcOutL0_240[2], gpcOutL0_189[0], gpcOutL0_188[1], gpcOutL0_187[2], gpcOutL0_133[0], gpcOutL0_132[1]}, gpcOutL1_54);
gpc006 gpcL1_55 ({gpcOutL0_190[0], gpcOutL0_189[1], gpcOutL0_188[2], gpcOutL0_134[0], gpcOutL0_133[1], gpcOutL0_132[2]}, gpcOutL1_55);
gpc006 gpcL1_56 ({gpcOutL0_191[0], gpcOutL0_190[1], gpcOutL0_189[2], gpcOutL0_135[0], gpcOutL0_134[1], gpcOutL0_133[2]}, gpcOutL1_56);
gpc006 gpcL1_57 ({gpcOutL0_229[0], gpcOutL0_191[1], gpcOutL0_190[2], gpcOutL0_136[0], gpcOutL0_135[1], gpcOutL0_134[2]}, gpcOutL1_57);
gpc006 gpcL1_58 ({gpcOutL0_241[0], gpcOutL0_229[1], gpcOutL0_191[2], gpcOutL0_137[0], gpcOutL0_136[1], gpcOutL0_135[2]}, gpcOutL1_58);
gpc006 gpcL1_59 ({gpcOutL0_253[0], gpcOutL0_241[1], gpcOutL0_229[2], gpcOutL0_138[0], gpcOutL0_137[1], gpcOutL0_136[2]}, gpcOutL1_59);
gpc006 gpcL1_60 ({gpcOutL0_253[1], gpcOutL0_242[0], gpcOutL0_241[2], gpcOutL0_139[0], gpcOutL0_138[1], gpcOutL0_137[2]}, gpcOutL1_60);
gpc006 gpcL1_61 ({gpcOutL0_242[1], gpcOutL0_140[0], gpcOutL0_139[1], gpcOutL0_138[2], gpcOutL0_68[0], gpcOutL0_67[1]}, gpcOutL1_61);
gpc006 gpcL1_62 ({gpcOutL0_242[2], gpcOutL0_141[0], gpcOutL0_140[1], gpcOutL0_139[2], gpcOutL0_69[0], gpcOutL0_68[1]}, gpcOutL1_62);
gpc006 gpcL1_63 ({gpcOutL0_142[0], gpcOutL0_141[1], gpcOutL0_140[2], gpcOutL0_70[0], gpcOutL0_69[1], gpcOutL0_68[2]}, gpcOutL1_63);
gpc006 gpcL1_64 ({gpcOutL0_143[0], gpcOutL0_142[1], gpcOutL0_141[2], gpcOutL0_71[0], gpcOutL0_70[1], gpcOutL0_69[2]}, gpcOutL1_64);
gpc006 gpcL1_65 ({gpcOutL0_230[0], gpcOutL0_143[1], gpcOutL0_142[2], gpcOutL0_72[0], gpcOutL0_71[1], gpcOutL0_70[2]}, gpcOutL1_65);
gpc006 gpcL1_66 ({gpcOutL0_243[0], gpcOutL0_230[1], gpcOutL0_143[2], gpcOutL0_73[0], gpcOutL0_72[1], gpcOutL0_71[2]}, gpcOutL1_66);
gpc006 gpcL1_67 ({gpcOutL0_254[0], gpcOutL0_243[1], gpcOutL0_230[2], gpcOutL0_74[0], gpcOutL0_73[1], gpcOutL0_72[2]}, gpcOutL1_67);
gpc006 gpcL1_68 ({gpcOutL0_254[1], gpcOutL0_244[0], gpcOutL0_243[2], gpcOutL0_75[0], gpcOutL0_74[1], gpcOutL0_73[2]}, gpcOutL1_68);
gpc006 gpcL1_69 ({gpcOutL0_244[2], gpcOutL0_77[0], gpcOutL0_76[1], gpcOutL0_75[2], pp223[3], pp215[5]}, gpcOutL1_69);
gpc006 gpcL1_70 ({gpcOutL0_94[0], gpcOutL0_93[1], gpcOutL0_92[2], gpcOutL0_22[0], gpcOutL0_21[1], gpcOutL0_20[2]}, gpcOutL1_70);
gpc006 gpcL1_71 ({gpcOutL0_94[1], gpcOutL0_93[2], gpcOutL0_23[0], gpcOutL0_22[1], gpcOutL0_21[2], pp7[3]}, gpcOutL1_71);
gpc006 gpcL1_72 ({gpcOutL0_96[0], gpcOutL0_95[1], gpcOutL0_94[2], gpcOutL0_24[0], gpcOutL0_23[1], gpcOutL0_22[2]}, gpcOutL1_72);
gpc006 gpcL1_73 ({gpcOutL0_98[0], gpcOutL0_97[1], gpcOutL0_96[2], gpcOutL0_26[0], gpcOutL0_25[1], gpcOutL0_24[2]}, gpcOutL1_73);
gpc006 gpcL1_74 ({gpcOutL0_99[0], gpcOutL0_98[1], gpcOutL0_97[2], gpcOutL0_27[0], gpcOutL0_26[1], gpcOutL0_25[2]}, gpcOutL1_74);
gpc006 gpcL1_75 ({gpcOutL0_100[0], gpcOutL0_99[1], gpcOutL0_98[2], gpcOutL0_28[0], gpcOutL0_27[1], gpcOutL0_26[2]}, gpcOutL1_75);
gpc006 gpcL1_76 ({gpcOutL0_101[0], gpcOutL0_100[1], gpcOutL0_99[2], gpcOutL0_29[0], gpcOutL0_28[1], gpcOutL0_27[2]}, gpcOutL1_76);
gpc006 gpcL1_77 ({gpcOutL0_102[0], gpcOutL0_101[1], gpcOutL0_100[2], gpcOutL0_30[0], gpcOutL0_29[1], gpcOutL0_28[2]}, gpcOutL1_77);
gpc006 gpcL1_78 ({gpcOutL0_103[0], gpcOutL0_102[1], gpcOutL0_101[2], gpcOutL0_31[0], gpcOutL0_30[1], gpcOutL0_29[2]}, gpcOutL1_78);
gpc006 gpcL1_79 ({gpcOutL0_104[0], gpcOutL0_103[1], gpcOutL0_102[2], gpcOutL0_32[0], gpcOutL0_31[1], gpcOutL0_30[2]}, gpcOutL1_79);
gpc006 gpcL1_80 ({gpcOutL0_105[0], gpcOutL0_104[1], gpcOutL0_103[2], gpcOutL0_33[0], gpcOutL0_32[1], gpcOutL0_31[2]}, gpcOutL1_80);
gpc006 gpcL1_81 ({gpcOutL0_106[0], gpcOutL0_105[1], gpcOutL0_104[2], gpcOutL0_34[0], gpcOutL0_33[1], gpcOutL0_32[2]}, gpcOutL1_81);
gpc006 gpcL1_82 ({gpcOutL0_107[0], gpcOutL0_106[1], gpcOutL0_105[2], gpcOutL0_35[0], gpcOutL0_34[1], gpcOutL0_33[2]}, gpcOutL1_82);
gpc006 gpcL1_83 ({gpcOutL0_108[0], gpcOutL0_107[1], gpcOutL0_106[2], gpcOutL0_36[0], gpcOutL0_35[1], gpcOutL0_34[2]}, gpcOutL1_83);
gpc006 gpcL1_84 ({gpcOutL0_109[0], gpcOutL0_108[1], gpcOutL0_107[2], gpcOutL0_37[0], gpcOutL0_36[1], gpcOutL0_35[2]}, gpcOutL1_84);
gpc006 gpcL1_85 ({gpcOutL0_110[0], gpcOutL0_109[1], gpcOutL0_108[2], gpcOutL0_38[0], gpcOutL0_37[1], gpcOutL0_36[2]}, gpcOutL1_85);
gpc006 gpcL1_86 ({gpcOutL0_111[0], gpcOutL0_110[1], gpcOutL0_109[2], gpcOutL0_39[0], gpcOutL0_38[1], gpcOutL0_37[2]}, gpcOutL1_86);
gpc006 gpcL1_87 ({gpcOutL0_112[0], gpcOutL0_111[1], gpcOutL0_110[2], gpcOutL0_40[0], gpcOutL0_39[1], gpcOutL0_38[2]}, gpcOutL1_87);
gpc006 gpcL1_88 ({gpcOutL0_113[0], gpcOutL0_112[1], gpcOutL0_111[2], gpcOutL0_41[0], gpcOutL0_40[1], gpcOutL0_39[2]}, gpcOutL1_88);
gpc006 gpcL1_89 ({gpcOutL0_114[0], gpcOutL0_113[1], gpcOutL0_112[2], gpcOutL0_42[0], gpcOutL0_41[1], gpcOutL0_40[2]}, gpcOutL1_89);
gpc006 gpcL1_90 ({gpcOutL0_115[0], gpcOutL0_114[1], gpcOutL0_113[2], gpcOutL0_43[0], gpcOutL0_42[1], gpcOutL0_41[2]}, gpcOutL1_90);
gpc006 gpcL1_91 ({gpcOutL0_116[0], gpcOutL0_115[1], gpcOutL0_114[2], gpcOutL0_44[0], gpcOutL0_43[1], gpcOutL0_42[2]}, gpcOutL1_91);
gpc006 gpcL1_92 ({gpcOutL0_117[0], gpcOutL0_116[1], gpcOutL0_115[2], gpcOutL0_45[0], gpcOutL0_44[1], gpcOutL0_43[2]}, gpcOutL1_92);
gpc006 gpcL1_93 ({gpcOutL0_118[0], gpcOutL0_117[1], gpcOutL0_116[2], gpcOutL0_46[0], gpcOutL0_45[1], gpcOutL0_44[2]}, gpcOutL1_93);
gpc006 gpcL1_94 ({gpcOutL0_119[0], gpcOutL0_118[1], gpcOutL0_117[2], gpcOutL0_47[0], gpcOutL0_46[1], gpcOutL0_45[2]}, gpcOutL1_94);
gpc006 gpcL1_95 ({gpcOutL0_120[0], gpcOutL0_119[1], gpcOutL0_118[2], gpcOutL0_48[0], gpcOutL0_47[1], gpcOutL0_46[2]}, gpcOutL1_95);
gpc006 gpcL1_96 ({gpcOutL0_121[0], gpcOutL0_120[1], gpcOutL0_119[2], gpcOutL0_49[0], gpcOutL0_48[1], gpcOutL0_47[2]}, gpcOutL1_96);
gpc006 gpcL1_97 ({gpcOutL0_122[0], gpcOutL0_121[1], gpcOutL0_120[2], gpcOutL0_50[0], gpcOutL0_49[1], gpcOutL0_48[2]}, gpcOutL1_97);
gpc006 gpcL1_98 ({gpcOutL0_123[0], gpcOutL0_122[1], gpcOutL0_121[2], gpcOutL0_51[0], gpcOutL0_50[1], gpcOutL0_49[2]}, gpcOutL1_98);
gpc006 gpcL1_99 ({gpcOutL0_124[0], gpcOutL0_123[1], gpcOutL0_122[2], gpcOutL0_52[0], gpcOutL0_51[1], gpcOutL0_50[2]}, gpcOutL1_99);
gpc006 gpcL1_100 ({gpcOutL0_125[0], gpcOutL0_124[1], gpcOutL0_123[2], gpcOutL0_53[0], gpcOutL0_52[1], gpcOutL0_51[2]}, gpcOutL1_100);
gpc006 gpcL1_101 ({gpcOutL0_126[0], gpcOutL0_125[1], gpcOutL0_124[2], gpcOutL0_54[0], gpcOutL0_53[1], gpcOutL0_52[2]}, gpcOutL1_101);
gpc006 gpcL1_102 ({gpcOutL0_127[0], gpcOutL0_126[1], gpcOutL0_125[2], gpcOutL0_55[0], gpcOutL0_54[1], gpcOutL0_53[2]}, gpcOutL1_102);
gpc006 gpcL1_103 ({gpcOutL0_128[0], gpcOutL0_127[1], gpcOutL0_126[2], gpcOutL0_56[0], gpcOutL0_55[1], gpcOutL0_54[2]}, gpcOutL1_103);
gpc006 gpcL1_104 ({gpcOutL0_129[0], gpcOutL0_128[1], gpcOutL0_127[2], gpcOutL0_57[0], gpcOutL0_56[1], gpcOutL0_55[2]}, gpcOutL1_104);
gpc006 gpcL1_105 ({gpcOutL0_130[0], gpcOutL0_129[1], gpcOutL0_128[2], gpcOutL0_58[0], gpcOutL0_57[1], gpcOutL0_56[2]}, gpcOutL1_105);
gpc006 gpcL1_106 ({gpcOutL0_131[0], gpcOutL0_130[1], gpcOutL0_129[2], gpcOutL0_59[0], gpcOutL0_58[1], gpcOutL0_57[2]}, gpcOutL1_106);
gpc006 gpcL1_107 ({gpcOutL0_131[2], gpcOutL0_61[0], gpcOutL0_60[1], gpcOutL0_59[2], pp159[3], pp151[5]}, gpcOutL1_107);
gpc015 gpcL1_108 ({gpcOutL0_248[0], gpcOutL0_256[2], gpcOutL0_234[0], gpcOutL0_4[0], gpcOutL0_3[1], gpcOutL0_2[2]}, gpcOutL1_108);
gpc015 gpcL1_109 ({gpcOutL0_92[1], gpcOutL0_91[1], gpcOutL0_90[2], gpcOutL0_20[0], gpcOutL0_19[1], gpcOutL0_18[2]}, gpcOutL1_109);
gpc005 gpcL1_110 ({gpcOutL0_235[0], gpcOutL0_225[1], gpcOutL0_7[0], gpcOutL0_6[1], gpcOutL0_5[2]}, gpcOutL1_110);
gpc005 gpcL1_111 ({gpcOutL0_96[1], gpcOutL0_95[2], gpcOutL0_25[0], gpcOutL0_24[1], gpcOutL0_23[2]}, gpcOutL1_111);
gpc005 gpcL1_112 ({gpcOutL0_130[2], gpcOutL0_60[0], gpcOutL0_59[1], gpcOutL0_58[2], pp151[4]}, gpcOutL1_112);
gpc005 gpcL1_113 ({gpcOutL0_244[1], gpcOutL0_76[0], gpcOutL0_75[1], gpcOutL0_74[2], pp215[4]}, gpcOutL1_113);
gpc014 gpcL1_114 ({gpcOutL0_256[0], gpcOutL0_233[2], gpcOutL0_1[0], gpcOutL0_0[1], pp1[5]}, gpcOutL1_114);
gpc014 gpcL1_115 ({gpcOutL0_88[2], gpcOutL0_17[0], gpcOutL0_16[1], gpcOutL0_15[2], pp5[5]}, gpcOutL1_115);
gpc014 gpcL1_116 ({gpcOutL0_63[0], gpcOutL0_62[0], gpcOutL0_61[1], gpcOutL0_60[2], pp159[4]}, gpcOutL1_116);
gpc014 gpcL1_117 ({gpcOutL0_79[0], gpcOutL0_78[0], gpcOutL0_77[1], gpcOutL0_76[2], pp223[4]}, gpcOutL1_117);
gpc023 gpcL1_118 ({gpcOutL0_256[1], gpcOutL0_3[0], gpcOutL0_2[0], gpcOutL0_1[1], gpcOutL0_0[2]}, gpcOutL1_118);
gpc023 gpcL1_119 ({gpcOutL0_14[1], gpcOutL0_13[2], gpcOutL0_14[0], gpcOutL0_13[1], gpcOutL0_12[2]}, gpcOutL1_119);
gpc023 gpcL1_120 ({gpcOutL0_89[2], gpcOutL0_19[0], gpcOutL0_18[0], gpcOutL0_17[1], gpcOutL0_16[2]}, gpcOutL1_120);
gpc023 gpcL1_121 ({gpcOutL0_64[0], gpcOutL0_63[1], gpcOutL0_62[1], gpcOutL0_61[2], pp159[5]}, gpcOutL1_121);
gpc023 gpcL1_122 ({gpcOutL0_66[0], gpcOutL0_65[1], gpcOutL0_65[0], gpcOutL0_64[1], gpcOutL0_63[2]}, gpcOutL1_122);
gpc023 gpcL1_123 ({gpcOutL0_66[2], pp183[4], gpcOutL0_67[0], gpcOutL0_66[1], gpcOutL0_65[2]}, gpcOutL1_123);
gpc023 gpcL1_124 ({gpcOutL0_231[0], gpcOutL0_79[1], gpcOutL0_78[1], gpcOutL0_77[2], pp223[5]}, gpcOutL1_124);
gpc023 gpcL1_125 ({gpcOutL0_255[0], gpcOutL0_245[1], gpcOutL0_245[0], gpcOutL0_231[1], gpcOutL0_79[2]}, gpcOutL1_125);
gpc023 gpcL1_126 ({gpcOutL0_246[1], pp247[4], gpcOutL0_255[1], gpcOutL0_246[0], gpcOutL0_245[2]}, gpcOutL1_126);
gpc003 gpcL1_127 ({gpcOutL0_234[1], gpcOutL0_5[0], gpcOutL0_4[1]}, gpcOutL1_127);
gpc003 gpcL1_128 ({gpcOutL0_16[0], gpcOutL0_15[1], gpcOutL0_14[2]}, gpcOutL1_128);
gpc003 gpcL1_129 ({gpcOutL0_91[2], gpcOutL0_21[0], gpcOutL0_20[1]}, gpcOutL1_129);
gpc003 gpcL1_130 ({gpcOutL0_67[2], pp191[3], pp183[5]}, gpcOutL1_130);
gpc003 gpcL1_131 ({gpcOutL0_246[2], pp255[3], pp247[5]}, gpcOutL1_131);
gpc022 gpcL1_132 ({gpcOutL0_12[1], gpcOutL0_11[2], gpcOutL0_11[1], gpcOutL0_10[2]}, gpcOutL1_132);
gpc222 gpcL1_133 ({gpcOutL0_247[1], gpcOutL0_232[2], gpcOutL0_247[0], gpcOutL0_232[1], gpcOutL0_259[2], gpcOutL0_232[0]}, gpcOutL1_133);

// level 2
wire [2:0]  gpcOutL2_0;
wire [2:0]  gpcOutL2_1;
wire [2:0]  gpcOutL2_2;
wire [2:0]  gpcOutL2_3;
wire [2:0]  gpcOutL2_4;
wire [2:0]  gpcOutL2_5;
wire [2:0]  gpcOutL2_6;
wire [2:0]  gpcOutL2_7;
wire [2:0]  gpcOutL2_8;
wire [2:0]  gpcOutL2_9;
wire [2:0]  gpcOutL2_10;
wire [2:0]  gpcOutL2_11;
wire [2:0]  gpcOutL2_12;
wire [2:0]  gpcOutL2_13;
wire [2:0]  gpcOutL2_14;
wire [2:0]  gpcOutL2_15;
wire [2:0]  gpcOutL2_16;
wire [2:0]  gpcOutL2_17;
wire [2:0]  gpcOutL2_18;
wire [2:0]  gpcOutL2_19;
wire [2:0]  gpcOutL2_20;
wire [2:0]  gpcOutL2_21;
wire [2:0]  gpcOutL2_22;
wire [2:0]  gpcOutL2_23;
wire [2:0]  gpcOutL2_24;
wire [2:0]  gpcOutL2_25;
wire [2:0]  gpcOutL2_26;
wire [2:0]  gpcOutL2_27;
wire [2:0]  gpcOutL2_28;
wire [2:0]  gpcOutL2_29;
wire [2:0]  gpcOutL2_30;
wire [2:0]  gpcOutL2_31;
wire [2:0]  gpcOutL2_32;
wire [2:0]  gpcOutL2_33;
wire [2:0]  gpcOutL2_34;
wire [2:0]  gpcOutL2_35;
wire [2:0]  gpcOutL2_36;
wire [2:0]  gpcOutL2_37;
wire [2:0]  gpcOutL2_38;
wire [2:0]  gpcOutL2_39;
wire [2:0]  gpcOutL2_40;
wire [2:0]  gpcOutL2_41;
wire [2:0]  gpcOutL2_42;
wire [2:0]  gpcOutL2_43;
wire [2:0]  gpcOutL2_44;
wire [2:0]  gpcOutL2_45;
wire [2:0]  gpcOutL2_46;
wire [2:0]  gpcOutL2_47;
wire [2:0]  gpcOutL2_48;
wire [2:0]  gpcOutL2_49;
wire [2:0]  gpcOutL2_50;
wire [2:0]  gpcOutL2_51;
wire [2:0]  gpcOutL2_52;
wire [2:0]  gpcOutL2_53;
wire [2:0]  gpcOutL2_54;
wire [2:0]  gpcOutL2_55;
wire [2:0]  gpcOutL2_56;
wire [2:0]  gpcOutL2_57;
wire [2:0]  gpcOutL2_58;
wire [2:0]  gpcOutL2_59;
wire [2:0]  gpcOutL2_60;
wire [2:0]  gpcOutL2_61;
wire [2:0]  gpcOutL2_62;
wire [1:0]  gpcOutL2_63;
wire [1:0]  gpcOutL2_64;
wire [1:0]  gpcOutL2_65;
wire [1:0]  gpcOutL2_66;
wire [1:0]  gpcOutL2_67;
wire [3:0]  gpcOutL2_68;

gpc006 gpcL2_0 ({gpcOutL1_120[1], gpcOutL1_115[2], gpcOutL1_12[0], gpcOutL1_11[1], gpcOutL1_10[2], gpcOutL0_18[1]}, gpcOutL2_0);
gpc006 gpcL2_1 ({gpcOutL1_129[0], gpcOutL1_109[1], gpcOutL1_14[0], gpcOutL1_13[1], gpcOutL1_12[2], gpcOutL0_19[2]}, gpcOutL2_1);
gpc006 gpcL2_2 ({gpcOutL1_129[1], gpcOutL1_109[2], gpcOutL1_70[0], gpcOutL1_15[0], gpcOutL1_14[1], gpcOutL1_13[2]}, gpcOutL2_2);
gpc006 gpcL2_3 ({gpcOutL1_72[0], gpcOutL1_71[1], gpcOutL1_70[2], gpcOutL1_17[0], gpcOutL1_16[1], gpcOutL1_15[2]}, gpcOutL2_3);
gpc006 gpcL2_4 ({gpcOutL1_111[0], gpcOutL1_72[1], gpcOutL1_71[2], gpcOutL1_18[0], gpcOutL1_17[1], gpcOutL1_16[2]}, gpcOutL2_4);
gpc006 gpcL2_5 ({gpcOutL1_111[1], gpcOutL1_73[0], gpcOutL1_72[2], gpcOutL1_19[0], gpcOutL1_18[1], gpcOutL1_17[2]}, gpcOutL2_5);
gpc006 gpcL2_6 ({gpcOutL1_111[2], gpcOutL1_74[0], gpcOutL1_73[1], gpcOutL1_20[0], gpcOutL1_19[1], gpcOutL1_18[2]}, gpcOutL2_6);
gpc006 gpcL2_7 ({gpcOutL1_75[0], gpcOutL1_74[1], gpcOutL1_73[2], gpcOutL1_21[0], gpcOutL1_20[1], gpcOutL1_19[2]}, gpcOutL2_7);
gpc006 gpcL2_8 ({gpcOutL1_76[0], gpcOutL1_75[1], gpcOutL1_74[2], gpcOutL1_22[0], gpcOutL1_21[1], gpcOutL1_20[2]}, gpcOutL2_8);
gpc006 gpcL2_9 ({gpcOutL1_77[0], gpcOutL1_76[1], gpcOutL1_75[2], gpcOutL1_23[0], gpcOutL1_22[1], gpcOutL1_21[2]}, gpcOutL2_9);
gpc006 gpcL2_10 ({gpcOutL1_78[0], gpcOutL1_77[1], gpcOutL1_76[2], gpcOutL1_24[0], gpcOutL1_23[1], gpcOutL1_22[2]}, gpcOutL2_10);
gpc006 gpcL2_11 ({gpcOutL1_79[0], gpcOutL1_78[1], gpcOutL1_77[2], gpcOutL1_25[0], gpcOutL1_24[1], gpcOutL1_23[2]}, gpcOutL2_11);
gpc006 gpcL2_12 ({gpcOutL1_80[0], gpcOutL1_79[1], gpcOutL1_78[2], gpcOutL1_26[0], gpcOutL1_25[1], gpcOutL1_24[2]}, gpcOutL2_12);
gpc006 gpcL2_13 ({gpcOutL1_81[0], gpcOutL1_80[1], gpcOutL1_79[2], gpcOutL1_27[0], gpcOutL1_26[1], gpcOutL1_25[2]}, gpcOutL2_13);
gpc006 gpcL2_14 ({gpcOutL1_82[0], gpcOutL1_81[1], gpcOutL1_80[2], gpcOutL1_28[0], gpcOutL1_27[1], gpcOutL1_26[2]}, gpcOutL2_14);
gpc006 gpcL2_15 ({gpcOutL1_83[0], gpcOutL1_82[1], gpcOutL1_81[2], gpcOutL1_29[0], gpcOutL1_28[1], gpcOutL1_27[2]}, gpcOutL2_15);
gpc006 gpcL2_16 ({gpcOutL1_84[0], gpcOutL1_83[1], gpcOutL1_82[2], gpcOutL1_30[0], gpcOutL1_29[1], gpcOutL1_28[2]}, gpcOutL2_16);
gpc006 gpcL2_17 ({gpcOutL1_85[0], gpcOutL1_84[1], gpcOutL1_83[2], gpcOutL1_31[0], gpcOutL1_30[1], gpcOutL1_29[2]}, gpcOutL2_17);
gpc006 gpcL2_18 ({gpcOutL1_86[0], gpcOutL1_85[1], gpcOutL1_84[2], gpcOutL1_32[0], gpcOutL1_31[1], gpcOutL1_30[2]}, gpcOutL2_18);
gpc006 gpcL2_19 ({gpcOutL1_87[0], gpcOutL1_86[1], gpcOutL1_85[2], gpcOutL1_33[0], gpcOutL1_32[1], gpcOutL1_31[2]}, gpcOutL2_19);
gpc006 gpcL2_20 ({gpcOutL1_88[0], gpcOutL1_87[1], gpcOutL1_86[2], gpcOutL1_34[0], gpcOutL1_33[1], gpcOutL1_32[2]}, gpcOutL2_20);
gpc006 gpcL2_21 ({gpcOutL1_89[0], gpcOutL1_88[1], gpcOutL1_87[2], gpcOutL1_35[0], gpcOutL1_34[1], gpcOutL1_33[2]}, gpcOutL2_21);
gpc006 gpcL2_22 ({gpcOutL1_90[0], gpcOutL1_89[1], gpcOutL1_88[2], gpcOutL1_36[0], gpcOutL1_35[1], gpcOutL1_34[2]}, gpcOutL2_22);
gpc006 gpcL2_23 ({gpcOutL1_91[0], gpcOutL1_90[1], gpcOutL1_89[2], gpcOutL1_37[0], gpcOutL1_36[1], gpcOutL1_35[2]}, gpcOutL2_23);
gpc006 gpcL2_24 ({gpcOutL1_92[0], gpcOutL1_91[1], gpcOutL1_90[2], gpcOutL1_38[0], gpcOutL1_37[1], gpcOutL1_36[2]}, gpcOutL2_24);
gpc006 gpcL2_25 ({gpcOutL1_93[0], gpcOutL1_92[1], gpcOutL1_91[2], gpcOutL1_39[0], gpcOutL1_38[1], gpcOutL1_37[2]}, gpcOutL2_25);
gpc006 gpcL2_26 ({gpcOutL1_94[0], gpcOutL1_93[1], gpcOutL1_92[2], gpcOutL1_40[0], gpcOutL1_39[1], gpcOutL1_38[2]}, gpcOutL2_26);
gpc006 gpcL2_27 ({gpcOutL1_95[0], gpcOutL1_94[1], gpcOutL1_93[2], gpcOutL1_41[0], gpcOutL1_40[1], gpcOutL1_39[2]}, gpcOutL2_27);
gpc006 gpcL2_28 ({gpcOutL1_96[0], gpcOutL1_95[1], gpcOutL1_94[2], gpcOutL1_42[0], gpcOutL1_41[1], gpcOutL1_40[2]}, gpcOutL2_28);
gpc006 gpcL2_29 ({gpcOutL1_97[0], gpcOutL1_96[1], gpcOutL1_95[2], gpcOutL1_43[0], gpcOutL1_42[1], gpcOutL1_41[2]}, gpcOutL2_29);
gpc006 gpcL2_30 ({gpcOutL1_98[0], gpcOutL1_97[1], gpcOutL1_96[2], gpcOutL1_44[0], gpcOutL1_43[1], gpcOutL1_42[2]}, gpcOutL2_30);
gpc006 gpcL2_31 ({gpcOutL1_99[0], gpcOutL1_98[1], gpcOutL1_97[2], gpcOutL1_45[0], gpcOutL1_44[1], gpcOutL1_43[2]}, gpcOutL2_31);
gpc006 gpcL2_32 ({gpcOutL1_100[0], gpcOutL1_99[1], gpcOutL1_98[2], gpcOutL1_46[0], gpcOutL1_45[1], gpcOutL1_44[2]}, gpcOutL2_32);
gpc006 gpcL2_33 ({gpcOutL1_101[0], gpcOutL1_100[1], gpcOutL1_99[2], gpcOutL1_47[0], gpcOutL1_46[1], gpcOutL1_45[2]}, gpcOutL2_33);
gpc006 gpcL2_34 ({gpcOutL1_102[0], gpcOutL1_101[1], gpcOutL1_100[2], gpcOutL1_48[0], gpcOutL1_47[1], gpcOutL1_46[2]}, gpcOutL2_34);
gpc006 gpcL2_35 ({gpcOutL1_103[0], gpcOutL1_102[1], gpcOutL1_101[2], gpcOutL1_49[0], gpcOutL1_48[1], gpcOutL1_47[2]}, gpcOutL2_35);
gpc006 gpcL2_36 ({gpcOutL1_104[0], gpcOutL1_103[1], gpcOutL1_102[2], gpcOutL1_50[0], gpcOutL1_49[1], gpcOutL1_48[2]}, gpcOutL2_36);
gpc006 gpcL2_37 ({gpcOutL1_105[0], gpcOutL1_104[1], gpcOutL1_103[2], gpcOutL1_51[0], gpcOutL1_50[1], gpcOutL1_49[2]}, gpcOutL2_37);
gpc006 gpcL2_38 ({gpcOutL1_106[0], gpcOutL1_105[1], gpcOutL1_104[2], gpcOutL1_52[0], gpcOutL1_51[1], gpcOutL1_50[2]}, gpcOutL2_38);
gpc006 gpcL2_39 ({gpcOutL1_112[0], gpcOutL1_106[1], gpcOutL1_105[2], gpcOutL1_53[0], gpcOutL1_52[1], gpcOutL1_51[2]}, gpcOutL2_39);
gpc006 gpcL2_40 ({gpcOutL1_112[1], gpcOutL1_107[0], gpcOutL1_106[2], gpcOutL1_54[0], gpcOutL1_53[1], gpcOutL1_52[2]}, gpcOutL2_40);
gpc006 gpcL2_41 ({gpcOutL1_116[0], gpcOutL1_112[2], gpcOutL1_107[1], gpcOutL1_55[0], gpcOutL1_54[1], gpcOutL1_53[2]}, gpcOutL2_41);
gpc006 gpcL2_42 ({gpcOutL1_121[0], gpcOutL1_116[1], gpcOutL1_107[2], gpcOutL1_56[0], gpcOutL1_55[1], gpcOutL1_54[2]}, gpcOutL2_42);
gpc006 gpcL2_43 ({gpcOutL1_121[1], gpcOutL1_116[2], gpcOutL1_57[0], gpcOutL1_56[1], gpcOutL1_55[2], gpcOutL0_62[2]}, gpcOutL2_43);
gpc015 gpcL2_44 ({gpcOutL1_119[1], gpcOutL1_132[2], gpcOutL1_119[0], gpcOutL1_7[0], gpcOutL1_6[1], gpcOutL1_5[2]}, gpcOutL2_44);
gpc015 gpcL2_45 ({gpcOutL1_128[1], gpcOutL1_128[0], gpcOutL1_119[2], gpcOutL1_9[0], gpcOutL1_8[1], gpcOutL1_7[2]}, gpcOutL2_45);
gpc015 gpcL2_46 ({gpcOutL0_17[2], gpcOutL1_120[0], gpcOutL1_115[1], gpcOutL1_11[0], gpcOutL1_10[1], gpcOutL1_9[2]}, gpcOutL2_46);
gpc015 gpcL2_47 ({gpcOutL1_122[1], gpcOutL1_122[0], gpcOutL1_121[2], gpcOutL1_58[0], gpcOutL1_57[1], gpcOutL1_56[2]}, gpcOutL2_47);
gpc015 gpcL2_48 ({gpcOutL1_123[1], gpcOutL1_123[0], gpcOutL1_122[2], gpcOutL1_60[0], gpcOutL1_59[1], gpcOutL1_58[2]}, gpcOutL2_48);
gpc015 gpcL2_49 ({gpcOutL1_130[1], gpcOutL1_130[0], gpcOutL1_123[2], gpcOutL1_62[0], gpcOutL1_61[1], gpcOutL1_60[2]}, gpcOutL2_49);
gpc005 gpcL2_50 ({gpcOutL1_120[2], gpcOutL1_109[0], gpcOutL1_13[0], gpcOutL1_12[1], gpcOutL1_11[2]}, gpcOutL2_50);
gpc005 gpcL2_51 ({gpcOutL1_71[0], gpcOutL1_70[1], gpcOutL1_16[0], gpcOutL1_15[1], gpcOutL1_14[2]}, gpcOutL2_51);
gpc014 gpcL2_52 ({gpcOutL1_118[2], gpcOutL1_118[1], gpcOutL1_114[2], gpcOutL0_2[1], gpcOutL0_1[2]}, gpcOutL2_52);
gpc014 gpcL2_53 ({gpcOutL1_3[0], gpcOutL1_110[2], gpcOutL1_2[0], gpcOutL1_1[1], pp3[5]}, gpcOutL2_53);
gpc014 gpcL2_54 ({gpcOutL1_132[0], gpcOutL1_4[0], gpcOutL1_3[1], gpcOutL1_2[2], gpcOutL0_9[2]}, gpcOutL2_54);
gpc014 gpcL2_55 ({gpcOutL1_64[0], gpcOutL1_63[0], gpcOutL1_62[1], gpcOutL1_61[2], pp191[4]}, gpcOutL2_55);
gpc023 gpcL2_56 ({gpcOutL1_127[1], gpcOutL1_108[2], gpcOutL1_127[0], gpcOutL1_108[1], gpcOutL0_3[2]}, gpcOutL2_56);
gpc023 gpcL2_57 ({gpcOutL1_132[1], gpcOutL1_6[0], gpcOutL1_5[0], gpcOutL1_4[1], gpcOutL1_3[2]}, gpcOutL2_57);
gpc023 gpcL2_58 ({gpcOutL1_65[0], gpcOutL1_64[1], gpcOutL1_63[1], gpcOutL1_62[2], pp191[5]}, gpcOutL2_58);
gpc023 gpcL2_59 ({gpcOutL1_67[0], gpcOutL1_66[1], gpcOutL1_66[0], gpcOutL1_65[1], gpcOutL1_64[2]}, gpcOutL2_59);
gpc023 gpcL2_60 ({gpcOutL1_113[0], gpcOutL1_68[1], gpcOutL1_68[0], gpcOutL1_67[1], gpcOutL1_66[2]}, gpcOutL2_60);
gpc023 gpcL2_61 ({gpcOutL1_117[0], gpcOutL1_113[2], gpcOutL1_113[1], gpcOutL1_69[0], gpcOutL1_68[2]}, gpcOutL2_61);
gpc023 gpcL2_62 ({gpcOutL1_124[1], gpcOutL1_117[2], gpcOutL1_124[0], gpcOutL1_117[1], gpcOutL1_69[2]}, gpcOutL2_62);
gpc003 gpcL2_63 ({gpcOutL1_2[1], gpcOutL1_1[2], gpcOutL0_8[2]}, gpcOutL2_63);
gpc003 gpcL2_64 ({gpcOutL1_8[0], gpcOutL1_7[1], gpcOutL1_6[2]}, gpcOutL2_64);
gpc003 gpcL2_65 ({gpcOutL1_115[0], gpcOutL1_10[0], gpcOutL1_9[1]}, gpcOutL2_65);
gpc003 gpcL2_66 ({gpcOutL1_59[0], gpcOutL1_58[1], gpcOutL1_57[2]}, gpcOutL2_66);
gpc003 gpcL2_67 ({gpcOutL1_61[0], gpcOutL1_60[1], gpcOutL1_59[2]}, gpcOutL2_67);
gpc132 gpcL2_68 ({gpcOutL0_233[1], gpcOutL1_133[3], gpcOutL0_233[0], gpcOutL0_224[1], gpcOutL1_133[2], gpcOutL0_224[0]}, gpcOutL2_68);

// level 3
wire [2:0]  gpcOutL3_0;
wire [2:0]  gpcOutL3_1;
wire [2:0]  gpcOutL3_2;

gpc014 gpcL3_0 ({gpcOutL2_57[2], gpcOutL2_57[1], gpcOutL2_54[2], gpcOutL1_5[1], gpcOutL1_4[2]}, gpcOutL3_0);
gpc014 gpcL3_1 ({gpcOutL2_66[1], gpcOutL2_66[0], gpcOutL2_47[1], gpcOutL2_43[2], gpcOutL0_64[2]}, gpcOutL3_1);
gpc023 gpcL3_2 ({gpcOutL2_68[3], gpcOutL1_114[0], gpcOutL2_68[2], gpcOutL0_224[2], gpcOutL0_0[0]}, gpcOutL3_2);

// final adder
wire [85:0]  adderIn0;
wire [85:0]  adderIn1;
wire [85:0]  adderIn2;
wire [86:0]  adderOut;

assign adderIn0 = {pp255[5], gpcOutL1_131[1], gpcOutL1_131[0], gpcOutL1_126[1], gpcOutL1_126[0], gpcOutL1_125[1], gpcOutL2_62[2], gpcOutL2_62[1], gpcOutL2_62[0], gpcOutL2_61[1], gpcOutL2_61[0], gpcOutL2_60[1], gpcOutL2_60[0], gpcOutL2_59[1], gpcOutL2_59[0], gpcOutL2_58[1], gpcOutL2_58[0], gpcOutL2_55[0], gpcOutL2_67[1], gpcOutL3_1[2], gpcOutL3_1[1], gpcOutL3_1[0], gpcOutL2_47[0], gpcOutL2_43[0], gpcOutL2_42[0], gpcOutL2_41[0], gpcOutL2_40[0], gpcOutL2_39[0], gpcOutL2_38[0], gpcOutL2_37[0], gpcOutL2_36[0], gpcOutL2_35[0], gpcOutL2_34[0], gpcOutL2_33[0], gpcOutL2_32[0], gpcOutL2_31[0], gpcOutL2_30[0], gpcOutL2_29[0], gpcOutL2_28[0], gpcOutL2_27[0], gpcOutL2_26[0], gpcOutL2_25[0], gpcOutL2_24[0], gpcOutL2_23[0], gpcOutL2_22[0], gpcOutL2_21[0], gpcOutL2_20[0], gpcOutL2_19[0], gpcOutL2_18[0], gpcOutL2_17[0], gpcOutL2_16[0], gpcOutL2_15[0], gpcOutL2_14[0], gpcOutL2_13[0], gpcOutL2_12[0], gpcOutL2_11[0], gpcOutL2_10[0], gpcOutL2_9[0], gpcOutL2_8[0], gpcOutL2_7[0], gpcOutL2_6[0], gpcOutL2_5[0], gpcOutL2_51[2], gpcOutL2_51[1], gpcOutL2_51[0], gpcOutL2_50[2], gpcOutL2_50[1], gpcOutL2_50[0], gpcOutL2_46[1], gpcOutL2_65[1], gpcOutL2_65[0], gpcOutL2_64[1], gpcOutL3_0[2], gpcOutL3_0[1], gpcOutL3_0[0], gpcOutL2_57[0], gpcOutL2_63[1], gpcOutL2_63[0], gpcOutL2_53[0], gpcOutL1_110[1], gpcOutL2_56[2], gpcOutL2_56[1], gpcOutL2_56[0], gpcOutL2_52[1], gpcOutL2_52[0], gpcOutL3_2[2]};
assign adderIn1 = {1'b0, pp255[4], gpcOutL1_126[2], 1'b0, gpcOutL1_125[2], gpcOutL0_231[2], gpcOutL1_125[0], gpcOutL0_78[2], gpcOutL2_61[2], gpcOutL1_69[1], gpcOutL2_60[2], gpcOutL1_67[2], gpcOutL2_59[2], gpcOutL1_65[2], gpcOutL2_58[2], gpcOutL2_55[2], gpcOutL2_55[1], gpcOutL2_49[1], gpcOutL2_49[0], gpcOutL2_67[0], gpcOutL2_48[0], 1'b0, gpcOutL2_43[1], gpcOutL2_42[1], gpcOutL2_41[1], gpcOutL2_40[1], gpcOutL2_39[1], gpcOutL2_38[1], gpcOutL2_37[1], gpcOutL2_36[1], gpcOutL2_35[1], gpcOutL2_34[1], gpcOutL2_33[1], gpcOutL2_32[1], gpcOutL2_31[1], gpcOutL2_30[1], gpcOutL2_29[1], gpcOutL2_28[1], gpcOutL2_27[1], gpcOutL2_26[1], gpcOutL2_25[1], gpcOutL2_24[1], gpcOutL2_23[1], gpcOutL2_22[1], gpcOutL2_21[1], gpcOutL2_20[1], gpcOutL2_19[1], gpcOutL2_18[1], gpcOutL2_17[1], gpcOutL2_16[1], gpcOutL2_15[1], gpcOutL2_14[1], gpcOutL2_13[1], gpcOutL2_12[1], gpcOutL2_11[1], gpcOutL2_10[1], gpcOutL2_9[1], gpcOutL2_8[1], gpcOutL2_7[1], gpcOutL2_6[1], gpcOutL2_5[1], gpcOutL2_4[1], gpcOutL2_4[0], gpcOutL2_3[0], gpcOutL2_2[1], gpcOutL2_2[0], gpcOutL2_1[0], gpcOutL2_46[2], gpcOutL2_0[0], gpcOutL2_46[0], gpcOutL2_45[1], gpcOutL2_45[0], gpcOutL2_64[0], gpcOutL2_44[0], 1'b0, gpcOutL2_54[1], gpcOutL2_54[0], gpcOutL2_53[1], 1'b0, gpcOutL1_1[0], gpcOutL1_110[0], gpcOutL1_0[0], gpcOutL2_52[2], gpcOutL1_108[0], 1'b0, gpcOutL1_118[0]};
assign adderIn2 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, gpcOutL1_124[2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, gpcOutL1_63[2], gpcOutL2_49[2], 1'b0, gpcOutL2_48[2], gpcOutL2_48[1], gpcOutL2_47[2], 1'b0, gpcOutL2_42[2], gpcOutL2_41[2], gpcOutL2_40[2], gpcOutL2_39[2], gpcOutL2_38[2], gpcOutL2_37[2], gpcOutL2_36[2], gpcOutL2_35[2], gpcOutL2_34[2], gpcOutL2_33[2], gpcOutL2_32[2], gpcOutL2_31[2], gpcOutL2_30[2], gpcOutL2_29[2], gpcOutL2_28[2], gpcOutL2_27[2], gpcOutL2_26[2], gpcOutL2_25[2], gpcOutL2_24[2], gpcOutL2_23[2], gpcOutL2_22[2], gpcOutL2_21[2], gpcOutL2_20[2], gpcOutL2_19[2], gpcOutL2_18[2], gpcOutL2_17[2], gpcOutL2_16[2], gpcOutL2_15[2], gpcOutL2_14[2], gpcOutL2_13[2], gpcOutL2_12[2], gpcOutL2_11[2], gpcOutL2_10[2], gpcOutL2_9[2], gpcOutL2_8[2], gpcOutL2_7[2], gpcOutL2_6[2], gpcOutL2_5[2], gpcOutL2_4[2], gpcOutL2_3[2], gpcOutL2_3[1], gpcOutL2_2[2], gpcOutL2_1[2], gpcOutL2_1[1], gpcOutL2_0[2], gpcOutL2_0[1], 1'b0, gpcOutL2_45[2], gpcOutL1_8[2], gpcOutL2_44[2], gpcOutL2_44[1], 1'b0, 1'b0, 1'b0, gpcOutL2_53[2], 1'b0, 1'b0, gpcOutL1_0[2], gpcOutL1_0[1], 1'b0, 1'b0, 1'b0, 1'b0, gpcOutL1_114[1]};
assign adderOut = adderIn0 + adderIn1 + adderIn2;

// multiplayer output
assign out = {adderOut[85:0], gpcOutL3_2[1], gpcOutL3_2[0], gpcOutL2_68[1], gpcOutL2_68[0], gpcOutL1_133[1], gpcOutL1_133[0], gpcOutL0_259[1], gpcOutL0_259[0], pp0[1], pp0[0]};

endmodule


/******************************************/

